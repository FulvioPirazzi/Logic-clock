//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "proj1 (copy).v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns


//: /symbolBegin: 3101448544
//: /iconBegin normal 365 5 14
//: /data "#define bitmap_width 29"
//: /data "#define bitmap_height 11"
//: /data "static unsigned char bitmap_bits[] = {"
//: /data "   0xff, 0x00, 0x00, 0x00, 0x02, 0x01, 0x00, 0x00, 0x02, 0x02, 0x00, 0x00,"
//: /data "   0x06, 0x04, 0x00, 0x00, 0x04, 0x04, 0x00, 0x00, 0x04, 0xfc, 0xff, 0x1f,"
//: /data "   0x04, 0x04, 0x00, 0x00, 0x04, 0x04, 0x00, 0x00, 0x06, 0x02, 0x00, 0x00,"
//: /data "   0x06, 0x01, 0x00, 0x00, 0xff, 0x00, 0x00, 0x00};"
//: /iconEnd
//: /iconBegin select 464 5 12
//: /data "#define bitmap_width 30"
//: /data "#define bitmap_height 15"
//: /data "static unsigned char bitmap_bits[] = {"
//: /data "   0x01, 0x00, 0x00, 0x00, 0xff, 0x00, 0x00, 0x00, 0x02, 0x03, 0x00, 0x00,"
//: /data "   0x02, 0x04, 0x00, 0x00, 0x04, 0x08, 0x00, 0x00, 0x74, 0x17, 0x00, 0x00,"
//: /data "   0x54, 0x15, 0x00, 0x00, 0x54, 0xf7, 0xff, 0x3f, 0x74, 0x19, 0x00, 0x00,"
//: /data "   0x04, 0x10, 0x00, 0x00, 0x04, 0x08, 0x00, 0x00, 0x02, 0x04, 0x00, 0x00,"
//: /data "   0x02, 0x03, 0x00, 0x00, 0xff, 0x00, 0x00, 0x00, 0x01, 0x00, 0x00, 0x00};"
//: /iconEnd
//: /port input A @(4, 14) /r:2
//: /port input B @(4, 24) /r:2
//: /port output Z @(34, 19) /r:0
//: /symbolEnd
//: /netlistBegin main
module main;    //: root_module
supply0 w4;    //: /sn:0 {0}(382,1722)(376,1722)(376,1687)(397,1687){1}
reg w104;    //: /sn:0 {0}(-812,638)(-817,638)(-817,600)(-169,600)(-169,-133)(254,-133)(254,-87){1}
reg w115;    //: /sn:0 {0}(301,-87)(301,-122)(-160,-122)(-160,604)(-921,604)(-921,922)(-548,922){1}
reg w117;    //: /sn:0 {0}(343,-87)(343,-127)(-165,-127)(-165,594)(-889,594)(-889,1860)(46,1860)(46,1841)(325,1841)(325,1867)(376,1867){1}
wire w32;    //: /sn:0 {0}(-6,802)(1,802)(1,793){1}
//: {2}(3,791)(37,791)(37,900)(-903,900)(-903,781)(-884,781){3}
//: {4}(1,789)(1,770)(112,770)(112,580){5}
//: {6}(112,576)(112,-227)(565,-227)(565,90){7}
//: {8}(563,92)(550,92){9}
//: {10}(565,94)(565,102){11}
//: {12}(567,104)(570,104)(570,114){13}
//: {14}(572,116)(575,116)(575,126){15}
//: {16}(573,128)(569,128)(569,128)(568,128){17}
//: {18}(577,128)(582,128)(582,138){19}
//: {20}(584,140)(587,140)(587,150){21}
//: {22}(589,152)(593,152)(593,164)(586,164){23}
//: {24}(585,152)(580,152){25}
//: {26}(580,140)(575,140)(575,140)(574,140){27}
//: {28}(568,116)(565,116)(565,116)(562,116){29}
//: {30}(563,104)(556,104){31}
//: {32}(110,578)(85,578)(85,578)(61,578){33}
wire w341;    //: /sn:0 {0}(32,1058)(17,1058){1}
//: {2}(15,1056)(15,940)(273,940)(273,828){3}
//: {4}(275,826)(305,826)(305,826)(547,826){5}
//: {6}(273,824)(273,670)(139,670)(139,-205)(1002,-205)(1002,-14)(796,-14)(796,-13){7}
//: {8}(794,-11)(792,-11){9}
//: {10}(796,-9)(796,0)(789,0){11}
//: {12}(785,0)(783,0)(783,0)(783,0){13}
//: {14}(787,2)(787,11)(781,11){15}
//: {16}(777,11)(774,11)(774,11)(774,11){17}
//: {18}(779,13)(779,22)(773,22){19}
//: {20}(769,22)(765,22)(765,22)(765,22){21}
//: {22}(771,24)(771,33)(763,33){23}
//: {24}(759,33)(756,33)(756,33)(756,33){25}
//: {26}(761,35)(761,44)(753,44){27}
//: {28}(749,44)(747,44)(747,44)(747,44){29}
//: {30}(1:751,46)(751,55)(744,55){31}
//: {32}(740,55)(738,55)(738,55)(738,55){33}
//: {34}(742,57)(742,66)(735,66){35}
//: {36}(731,66)(729,66)(729,66)(729,66){37}
//: {38}(733,68)(733,77)(729,77){39}
//: {40}(725,77)(721,77)(721,77)(720,77){41}
//: {42}(727,79)(727,88)(718,88){43}
//: {44}(714,88)(711,88)(711,88)(711,88){45}
//: {46}(716,90)(716,98)(702,98){47}
//: {48}(13,1058)(6,1058){49}
wire w364;    //: /sn:0 {0}(-115,1222)(-122,1222){1}
wire w270;    //: /sn:0 {0}(1121,2262)(1116,2262){1}
wire w160;    //: /sn:0 {0}(225,1061)(216,1061){1}
//: {2}(214,1059)(214,952)(279,952)(279,858){3}
//: {4}(281,856)(317,856)(317,856)(547,856){5}
//: {6}(279,854)(279,664)(145,664)(145,-199)(996,-199)(996,99)(846,99){7}
//: {8}(844,97)(844,88){9}
//: {10}(844,101)(844,103)(834,103){11}
//: {12}(832,101)(832,96)(832,96)(832,94){13}
//: {14}(832,105)(832,108)(822,108){15}
//: {16}(820,106)(820,103)(820,103)(820,100){17}
//: {18}(820,110)(820,113)(810,113){19}
//: {20}(808,111)(808,107)(808,107)(808,106){21}
//: {22}(808,115)(808,120)(798,120){23}
//: {24}(796,118)(796,112){25}
//: {26}(796,122)(796,127)(786,127){27}
//: {28}(784,125)(784,120)(784,120)(784,118){29}
//: {30}(784,129)(784,132)(774,132){31}
//: {32}(772,130)(772,127)(772,127)(772,124){33}
//: {34}(772,134)(772,137)(762,137){35}
//: {36}(760,135)(760,131)(760,131)(760,130){37}
//: {38}(760,139)(760,144)(750,144){39}
//: {40}(748,142)(748,137)(748,137)(748,136){41}
//: {42}(748,146)(748,149)(738,149){43}
//: {44}(736,147)(736,142){45}
//: {46}(736,151)(736,154)(724,154)(724,148){47}
//: {48}(212,1061)(204,1061){49}
wire w96;    //: /sn:0 {0}(1201,2240)(1192,2240){1}
//: {2}(1190,2238)(1190,2211)(1374,2211)(1374,1346){3}
//: {4}(1374,1342)(1374,550)(225,550)(225,-176)(559,-176)(559,-72)(554,-72){5}
//: {6}(1372,1344)(1197,1344){7}
//: {8}(1188,2240)(1180,2240){9}
wire [59:0] w45;    //: /sn:0 {0}(-94,540)(-105,540)(-105,721)(1302,721)(1302,1042)(1179,1042)(1179,1059)(#:1191,1059){1}
wire w73;    //: /sn:0 {0}(1197,944)(1282,944){1}
//: {2}(1284,942)(1284,645)(1037,645)(1037,299)(874,299)(874,290){3}
//: {4}(1284,946)(1284,1745)(929,1745)(929,1795){5}
//: {6}(931,1797)(942,1797){7}
//: {8}(927,1797)(919,1797){9}
wire w339;    //: /sn:0 {0}(98,1059)(86,1059){1}
//: {2}(84,1057)(84,945)(275,945)(275,838){3}
//: {4}(277,836)(310,836)(310,836)(547,836){5}
//: {6}(275,834)(275,668)(141,668)(141,-203)(1000,-203)(1000,26)(816,26){7}
//: {8}(814,24)(814,20){9}
//: {10}(814,28)(814,35)(806,35){11}
//: {12}(804,33)(804,30){13}
//: {14}(804,37)(804,44)(796,44){15}
//: {16}(794,42)(794,40){17}
//: {18}(794,46)(794,55)(785,55){19}
//: {20}(783,53)(783,49){21}
//: {22}(783,57)(783,63)(774,63){23}
//: {24}(772,61)(772,58){25}
//: {26}(772,65)(772,73)(764,73){27}
//: {28}(762,71)(762,69){29}
//: {30}(762,75)(762,82)(753,82){31}
//: {32}(751,80)(751,78){33}
//: {34}(751,84)(751,92)(742,92){35}
//: {36}(740,90)(740,88){37}
//: {38}(740,94)(740,101)(731,101){39}
//: {40}(729,99)(729,97){41}
//: {42}(729,103)(729,110)(720,110){43}
//: {44}(718,108)(718,107){45}
//: {46}(718,112)(718,118)(707,118)(707,116){47}
//: {48}(82,1059)(74,1059){49}
wire w359;    //: /sn:0 {0}(-377,1512)(-384,1512){1}
wire w320;    //: /sn:0 {0}(-248,1367)(-253,1367){1}
wire w16;    //: /sn:0 {0}(-791,641)(-785,641)(-785,848)(-774,848){1}
//: {2}(-770,848)(-712,848){3}
//: {4}(-708,848)(-647,848){5}
//: {6}(-643,848)(-636,848)(-636,848)(-580,848){7}
//: {8}(-576,848)(-547,848)(-547,848)(-513,848){9}
//: {10}(-509,848)(-451,848){11}
//: {12}(-447,848)(-386,848){13}
//: {14}(-382,848)(-321,848){15}
//: {16}(-317,848)(-310,848)(-310,848)(-254,848){17}
//: {18}(-250,848)(-218,848)(-218,848)(-187,848){19}
//: {20}(-183,848)(-137,848)(-137,848)(-125,848){21}
//: {22}(-121,848)(-57,848)(-57,825)(-48,825){23}
//: {24}(-123,846)(-123,824)(-111,824){25}
//: {26}(-185,846)(-185,823)(-175,823){27}
//: {28}(-252,846)(-252,822)(-241,822){29}
//: {30}(-319,846)(-319,821)(-309,821){31}
//: {32}(-384,846)(-384,820)(-374,820){33}
//: {34}(-449,846)(-449,819)(-437,819){35}
//: {36}(-511,846)(-511,818)(-501,818){37}
//: {38}(-578,846)(-578,817)(-567,817){39}
//: {40}(-645,846)(-645,816)(-635,816){41}
//: {42}(-710,846)(-710,815)(-698,815){43}
//: {44}(-772,846)(-772,814)(-762,814){45}
wire w56;    //: /sn:0 {0}(683,1940)(674,1940){1}
//: {2}(672,1938)(672,1869)(1304,1869)(1304,1026){3}
//: {4}(1304,1022)(1304,623)(682,623)(682,472)(698,472){5}
//: {6}(1302,1024)(1197,1024){7}
//: {8}(670,1940)(657,1940){9}
wire w218;    //: /sn:0 {0}(664,1963)(657,1963){1}
wire w81;    //: /sn:0 {0}(1244,2096)(1256,2096){1}
//: {2}(1258,2094)(1258,2062)(1349,2062)(1349,1236){3}
//: {4}(1349,1232)(1349,577)(234,577)(234,132)(323,132)(323,140){5}
//: {6}(1347,1234)(1197,1234){7}
//: {8}(1258,2098)(1258,2148)(477,2148)(477,2229)(487,2229){9}
wire w89;    //: /sn:0 {0}(547,896)(401,896)(401,896)(295,896){1}
//: {2}(293,894)(293,651)(153,651)(153,-191)(988,-191)(988,199)(864,199)(864,193){3}
//: {4}(864,189)(864,188){5}
//: {6}(862,191)(858,191)(858,192)(854,192){7}
//: {8}(852,190)(852,189){9}
//: {10}(850,192)(845,192)(845,193)(841,193){11}
//: {12}(839,191)(839,188)(839,188)(839,190){13}
//: {14}(837,193)(832,193)(832,194)(828,194){15}
//: {16}(826,192)(826,191)(826,191)(826,191){17}
//: {18}(824,194)(819,194)(819,195)(815,195){19}
//: {20}(813,193)(813,192){21}
//: {22}(811,195)(807,195)(807,196)(803,196){23}
//: {24}(801,194)(801,193)(801,193)(801,193){25}
//: {26}(799,196)(794,196)(794,197)(790,197){27}
//: {28}(788,195)(788,194)(788,194)(788,194){29}
//: {30}(786,197)(782,197)(782,198)(778,198){31}
//: {32}(776,196)(776,195)(776,195)(776,195){33}
//: {34}(774,198)(770,198)(770,199)(766,199){35}
//: {36}(764,197)(764,196)(764,196)(764,196){37}
//: {38}(762,199)(757,199)(757,200)(753,200){39}
//: {40}(751,198)(751,197){41}
//: {42}(749,200)(738,200)(738,198){43}
//: {44}(293,898)(293,1137)(-307,1137)(-307,1194){45}
//: {46}(-305,1196)(-294,1196){47}
//: {48}(-309,1196)(-320,1196){49}
wire w387;    //: /sn:0 {0}(13,1081)(6,1081){1}
wire w19;    //: /sn:0 {0}(61,658)(83,658)(83,658)(94,658){1}
//: {2}(96,656)(96,-237)(1066,-237)(1066,221)(727,221){3}
//: {4}(725,219)(725,211){5}
//: {6}(723,221)(715,221){7}
//: {8}(713,219)(713,212)(713,212)(713,211){9}
//: {10}(711,221)(702,221){11}
//: {12}(700,219)(700,211){13}
//: {14}(698,221)(690,221){15}
//: {16}(688,219)(688,212)(688,212)(688,211){17}
//: {18}(686,221)(678,221){19}
//: {20}(676,219)(676,211){21}
//: {22}(674,221)(665,221){23}
//: {24}(663,219)(663,211){25}
//: {26}(661,221)(650,221)(650,211){27}
//: {28}(96,660)(96,746)(-514,746)(-514,792){29}
//: {30}(-512,794)(-501,794){31}
//: {32}(-516,794)(-525,794){33}
wire w183;    //: /sn:0 {0}(-426,1341)(-433,1341){1}
//: {2}(-435,1339)(-435,1266)(317,1266)(317,998){3}
//: {4}(319,996)(413,996)(413,996)(547,996){5}
//: {6}(317,994)(317,677)(744,677)(744,440){7}
//: {8}(746,438)(749,438)(749,438)(750,438){9}
//: {10}(742,438)(736,438)(736,429){11}
//: {12}(738,427)(740,427)(740,427)(742,427){13}
//: {14}(734,427)(728,427)(728,418){15}
//: {16}(730,416)(732,416)(732,416)(734,416){17}
//: {18}(726,416)(719,416)(719,406){19}
//: {20}(721,404)(728,404)(728,404)(727,404){21}
//: {22}(717,404)(710,404)(710,394){23}
//: {24}(712,392)(718,392)(718,392)(719,392){25}
//: {26}(708,392)(704,392)(704,383){27}
//: {28}(706,381)(711,381)(711,381)(711,381){29}
//: {30}(702,381)(697,381)(697,371){31}
//: {32}(699,369)(703,369)(703,369)(703,369){33}
//: {34}(695,369)(691,369)(691,359){35}
//: {36}(693,357)(696,357)(696,357)(695,357){37}
//: {38}(689,357)(684,357)(684,347){39}
//: {40}(686,345)(688,345)(688,345)(688,345){41}
//: {42}(682,345)(675,345)(675,335){43}
//: {44}(677,333)(679,333)(679,333)(680,333){45}
//: {46}(673,333)(670,333)(670,321)(673,321){47}
//: {48}(-437,1341)(-448,1341){49}
wire w376;    //: /sn:0 {0}(78,1372)(73,1372){1}
wire w151;    //: /sn:0 {0}(-228,1054)(-237,1054){1}
//: {2}(-239,1052)(-239,925)(265,925)(265,788){3}
//: {4}(267,786)(318,786)(318,786)(547,786){5}
//: {6}(265,784)(265,678)(131,678)(131,-213)(699,-213)(699,-68)(686,-68)(686,-58){7}
//: {8}(684,-56)(683,-56){9}
//: {10}(686,-54)(686,-50)(682,-50)(682,-46){11}
//: {12}(680,-44)(675,-44)(675,-44)(679,-44){13}
//: {14}(682,-42)(682,-37)(679,-37)(679,-33){15}
//: {16}(677,-31)(672,-31)(672,-31)(676,-31){17}
//: {18}(679,-29)(679,-24)(676,-24)(676,-20){19}
//: {20}(674,-18)(667,-18)(667,-18)(671,-18){21}
//: {22}(676,-16)(676,-7)(672,-7)(672,-7){23}
//: {24}(670,-5)(663,-5)(663,-5)(667,-5){25}
//: {26}(672,-3)(672,1)(669,1)(669,6){27}
//: {28}(667,8)(660,8)(660,8)(664,8){29}
//: {30}(669,10)(669,15)(666,15)(666,19){31}
//: {32}(664,21)(657,21)(657,21)(661,21){33}
//: {34}(666,23)(666,27)(663,27)(663,31){35}
//: {36}(661,33)(654,33)(654,33)(658,33){37}
//: {38}(663,35)(663,39)(658,39)(658,43){39}
//: {40}(656,45)(649,45)(649,45)(653,45){41}
//: {42}(658,47)(658,52)(654,52)(654,56){43}
//: {44}(652,58)(645,58)(645,58)(649,58){45}
//: {46}(654,60)(654,71)(646,71){47}
//: {48}(-241,1054)(-252,1054){49}
wire w383;    //: /sn:0 {0}(-313,1076)(-320,1076){1}
wire w0;    //: /sn:0 {0}(-295,1490)(-304,1490){1}
//: {2}(-306,1488)(-306,1420)(349,1420)(349,1138){3}
//: {4}(351,1136)(429,1136)(429,1136)(547,1136){5}
//: {6}(349,1134)(349,605)(273,605)(273,380)(386,380){7}
//: {8}(388,378)(388,371)(396,371){9}
//: {10}(398,373)(398,376){11}
//: {12}(398,369)(398,362)(406,362){13}
//: {14}(408,364)(408,366){15}
//: {16}(408,360)(408,351)(417,351){17}
//: {18}(419,353)(419,357){19}
//: {20}(419,349)(419,343)(428,343){21}
//: {22}(430,345)(430,348){23}
//: {24}(430,341)(430,333)(438,333){25}
//: {26}(440,335)(440,337){27}
//: {28}(440,331)(440,324)(449,324){29}
//: {30}(451,326)(451,328){31}
//: {32}(451,322)(451,314)(460,314){33}
//: {34}(462,316)(462,318){35}
//: {36}(462,312)(462,305)(471,305){37}
//: {38}(473,307)(473,309){39}
//: {40}(473,303)(473,296)(482,296){41}
//: {42}(484,298)(484,299){43}
//: {44}(484,294)(484,288)(495,288)(495,290){45}
//: {46}(388,382)(388,386){47}
//: {48}(-308,1490)(-321,1490){49}
wire w120;    //: /sn:0 {0}(427,0)(430,0){1}
//: {2}(432,-2)(432,-10)(425,-10){3}
//: {4}(423,-12)(423,-147)(184,-147)(184,619)(384,619)(384,1284){5}
//: {6}(386,1286)(446,1286)(446,1286)(547,1286){7}
//: {8}(384,1288)(384,1589)(-113,1589)(-113,1636){9}
//: {10}(-111,1638)(-103,1638){11}
//: {12}(-115,1638)(-124,1638){13}
//: {14}(421,-10)(417,-10){15}
//: {16}(434,0)(441,0)(441,8){17}
//: {18}(439,10)(437,10){19}
//: {20}(443,10)(452,10)(452,19){21}
//: {22}(450,21)(446,21){23}
//: {24}(454,21)(460,21)(460,30){25}
//: {26}(458,32)(455,32){27}
//: {28}(462,32)(470,32)(470,40){29}
//: {30}(468,42)(466,42){31}
//: {32}(472,42)(479,42)(479,51){33}
//: {34}(477,53)(475,53){35}
//: {36}(481,53)(489,53)(489,62){37}
//: {38}(487,64)(485,64){39}
//: {40}(491,64)(498,64)(498,73){41}
//: {42}(496,75)(494,75){43}
//: {44}(500,75)(507,75)(507,84){45}
//: {46}(505,86)(504,86){47}
//: {48}(509,86)(515,86)(515,97)(513,97){49}
wire w233;    //: /sn:0 {0}(4,1640)(18,1640){1}
//: {2}(22,1640)(30,1640){3}
//: {4}(20,1638)(20,1600)(388,1600)(388,1308){5}
//: {6}(390,1306)(448,1306)(448,1306)(547,1306){7}
//: {8}(388,1304)(388,615)(190,615)(190,-151)(495,-151)(495,-42){9}
//: {10}(497,-40)(499,-40)(499,-30){11}
//: {12}(497,-28)(492,-28)(492,-28)(490,-28){13}
//: {14}(501,-28)(504,-28)(504,-18){15}
//: {16}(502,-16)(499,-16)(499,-16)(496,-16){17}
//: {18}(506,-16)(509,-16)(509,-6){19}
//: {20}(507,-4)(503,-4)(503,-4)(502,-4){21}
//: {22}(511,-4)(516,-4)(516,6){23}
//: {24}(514,8)(508,8){25}
//: {26}(518,8)(523,8)(523,18){27}
//: {28}(521,20)(516,20)(516,20)(514,20){29}
//: {30}(525,20)(528,20)(528,30){31}
//: {32}(526,32)(523,32)(523,32)(520,32){33}
//: {34}(530,32)(533,32)(533,42){35}
//: {36}(531,44)(527,44)(527,44)(526,44){37}
//: {38}(535,44)(540,44)(540,54){39}
//: {40}(538,56)(533,56)(533,56)(532,56){41}
//: {42}(542,56)(545,56)(545,66){43}
//: {44}(543,68)(538,68){45}
//: {46}(547,68)(551,68)(551,80)(544,80){47}
//: {48}(493,-40)(484,-40){49}
wire w313;    //: /sn:0 {0}(11,1663)(4,1663){1}
wire w111;    //: /sn:0 {0}(547,886)(400,886)(400,886)(293,886){1}
//: {2}(291,884)(291,653)(151,653)(151,-193)(990,-193)(990,175)(862,175)(862,167){3}
//: {4}(862,163)(862,162)(862,162)(862,161){5}
//: {6}(860,165)(858,165)(858,166)(852,166){7}
//: {8}(850,164)(850,163){9}
//: {10}(848,166)(843,166)(843,168)(839,168){11}
//: {12}(837,166)(837,163)(837,163)(837,165){13}
//: {14}(835,168)(830,168)(830,171)(826,171){15}
//: {16}(824,169)(824,168)(824,168)(824,168){17}
//: {18}(822,171)(818,171)(818,174)(813,174){19}
//: {20}(811,172)(811,171){21}
//: {22}(809,174)(805,174)(805,176)(801,176){23}
//: {24}(799,174)(799,174)(799,174)(799,173){25}
//: {26}(797,176)(792,176)(792,178)(788,178){27}
//: {28}(786,176)(786,175)(786,175)(786,175){29}
//: {30}(784,178)(780,178)(780,181)(775,181){31}
//: {32}(773,179)(773,178)(773,178)(773,178){33}
//: {34}(771,181)(767,181)(767,183)(763,183){35}
//: {36}(761,181)(761,180)(761,180)(761,180){37}
//: {38}(759,183)(754,183)(754,185)(750,185){39}
//: {40}(748,183)(748,182){41}
//: {42}(748,187)(748,190)(735,190)(735,185){43}
//: {44}(291,888)(291,1133)(-370,1133)(-370,1193){45}
//: {46}(-368,1195)(-362,1195){47}
//: {48}(-372,1195)(-383,1195){49}
wire w171;    //: /sn:0 {0}(-164,1198)(-173,1198){1}
//: {2}(-175,1196)(-175,1146)(297,1146)(297,918){3}
//: {4}(299,916)(403,916)(403,916)(547,916){5}
//: {6}(297,914)(297,698)(976,698)(976,254)(862,254)(862,244){7}
//: {8}(862,240)(862,237){9}
//: {10}(860,242)(856,242)(856,240)(852,240){11}
//: {12}(850,238)(850,231)(850,231)(850,235){13}
//: {14}(848,240)(843,240)(843,239)(839,239){15}
//: {16}(837,237)(837,230)(837,230)(837,234){17}
//: {18}(835,239)(830,239)(830,237)(826,237){19}
//: {20}(824,235)(824,228)(824,228)(824,232){21}
//: {22}(822,237)(813,237)(813,236)(813,236){23}
//: {24}(811,234)(811,227)(811,227)(811,231){25}
//: {26}(809,236)(805,236)(805,235)(800,235){27}
//: {28}(798,233)(798,226)(798,226)(798,230){29}
//: {30}(796,235)(791,235)(791,234)(787,234){31}
//: {32}(785,232)(785,225)(785,225)(785,229){33}
//: {34}(783,234)(779,234)(779,233)(775,233){35}
//: {36}(773,231)(773,224)(773,224)(773,228){37}
//: {38}(771,233)(767,233)(767,232)(763,232){39}
//: {40}(761,230)(761,223)(761,223)(761,227){41}
//: {42}(759,232)(754,232)(754,230)(750,230){43}
//: {44}(748,228)(748,225){45}
//: {46}(746,230)(738,230)(738,230)(735,230)(735,224){47}
//: {48}(-177,1198)(-186,1198){49}
wire w368;    //: /sn:0 {0}(-52,1080)(-59,1080){1}
wire w168;    //: /sn:0 {0}(602,1815)(595,1815){1}
wire w287;    //: /sn:0 {0}(162,1203)(154,1203){1}
//: {2}(152,1201)(152,1167)(307,1167)(307,968){3}
//: {4}(309,966)(408,966)(408,966)(547,966){5}
//: {6}(307,964)(307,688)(986,688)(986,374)(832,374){7}
//: {8}(830,372)(830,369){9}
//: {10}(828,374)(818,374)(818,369){11}
//: {12}(818,365)(818,362){13}
//: {14}(816,367)(806,367)(806,362){15}
//: {16}(806,358)(806,354){17}
//: {18}(804,360)(794,360)(794,355){19}
//: {20}(794,351)(794,347){21}
//: {22}(792,353)(782,353)(782,348){23}
//: {24}(782,344)(782,340)(782,340)(782,339){25}
//: {26}(780,346)(770,346)(770,339){27}
//: {28}(770,335)(770,331)(770,331)(770,331){29}
//: {30}(768,337)(1:758,337)(758,332){31}
//: {32}(758,328)(758,323){33}
//: {34}(756,330)(746,330)(746,323){35}
//: {36}(746,319)(746,315)(746,315)(746,315){37}
//: {38}(744,321)(734,321)(734,315){39}
//: {40}(734,311)(734,308)(734,308)(734,308){41}
//: {42}(732,313)(723,313)(723,308){43}
//: {44}(723,304)(723,299)(723,299)(723,299){45}
//: {46}(721,306)(714,306)(714,292){47}
//: {48}(150,1203)(140,1203){49}
wire w237;    //: /sn:0 {0}(862,2113)(855,2113){1}
wire w119;    //: /sn:0 {0}(1243,2241)(1259,2241)(1259,2230){1}
//: {2}(1261,2228)(1276,2228)(1276,2310)(273,2310)(273,1823){3}
//: {4}(1259,2226)(1259,2215)(1376,2215)(1376,1356){5}
//: {6}(1376,1352)(1376,548)(227,548)(227,-178)(585,-178)(585,-72)(582,-72){7}
//: {8}(1374,1354)(1197,1354){9}
wire w54;    //: /sn:0 {0}(552,1938)(545,1938){1}
//: {2}(543,1936)(543,1862)(1300,1862)(1300,1006){3}
//: {4}(1300,1002)(1300,627)(739,627)(739,451)(758,451){5}
//: {6}(1298,1004)(1197,1004){7}
//: {8}(541,1938)(530,1938){9}
wire w327;    //: /sn:0 {0}(-115,1079)(-122,1079){1}
wire w67;    //: /sn:0 {0}(-48,801)(-57,801){1}
//: {2}(-59,799)(-59,767)(110,767)(110,590){3}
//: {4}(110,586)(110,128)(490,128){5}
//: {6}(494,128)(504,128)(504,132){7}
//: {8}(506,134)(516,134)(516,137){9}
//: {10}(516,141)(516,150){11}
//: {12}(518,139)(528,139)(528,143){13}
//: {14}(528,147)(528,156){15}
//: {16}(530,145)(540,145)(540,149){17}
//: {18}(540,153)(540,162){19}
//: {20}(542,151)(552,151)(552,157){21}
//: {22}(554,159)(564,159)(564,174){23}
//: {24}(552,161)(552,168){25}
//: {26}(504,136)(504,140)(504,140)(504,144){27}
//: {28}(492,130)(492,138){29}
//: {30}(108,588)(95,588)(95,588)(61,588){31}
//: {32}(-61,801)(-69,801){33}
wire w90;    //: /sn:0 {0}(917,2236)(925,2236){1}
//: {2}(929,2236)(940,2236){3}
//: {4}(927,2234)(927,2191)(1366,2191)(1366,1306){5}
//: {6}(1366,1302)(1366,558)(217,558)(217,-168)(449,-168)(449,-42)(441,-42){7}
//: {8}(1364,1304)(1197,1304){9}
wire w294;    //: /sn:0 {0}(-247,1077)(-252,1077){1}
wire w176;    //: /sn:0 {0}(665,1816)(658,1816){1}
wire w174;    //: /sn:0 {0}(547,936)(405,936)(405,936)(303,936){1}
//: {2}(301,934)(301,694)(980,694)(980,294)(860,294)(860,292){3}
//: {4}(860,288)(860,287){5}
//: {6}(858,290)(854,290)(854,286)(850,286){7}
//: {8}(848,284)(848,279)(848,279)(848,283){9}
//: {10}(846,286)(841,286)(841,283)(837,283){11}
//: {12}(835,281)(835,276)(835,276)(835,280){13}
//: {14}(833,283)(828,283)(828,280)(824,280){15}
//: {16}(822,278)(822,271)(822,271)(822,275){17}
//: {18}(820,280)(811,280)(811,276)(811,276){19}
//: {20}(809,274)(809,267)(809,267)(809,271){21}
//: {22}(807,276)(803,276)(803,273)(798,273){23}
//: {24}(796,271)(796,264)(796,264)(796,268){25}
//: {26}(794,273)(789,273)(789,270)(785,270){27}
//: {28}(783,268)(783,261)(783,261)(783,265){29}
//: {30}(781,270)(777,270)(777,267)(773,267){31}
//: {32}(771,265)(771,258)(771,258)(771,262){33}
//: {34}(769,267)(765,267)(765,262)(761,262){35}
//: {36}(759,260)(759,253)(759,253)(759,257){37}
//: {38}(757,262)(752,262)(752,258)(748,258){39}
//: {40}(746,256)(746,249)(746,249)(746,253){41}
//: {42}(744,258)(733,258)(733,250){43}
//: {44}(301,938)(301,1154)(-49,1154)(-49,1198){45}
//: {46}(-47,1200)(-36,1200){47}
//: {48}(-51,1200)(-59,1200){49}
wire w20;    //: /sn:0 {0}(-720,791)(-712,791){1}
//: {2}(-708,791)(-698,791){3}
//: {4}(-710,789)(-710,737)(90,737)(90,690){5}
//: {6}(90,686)(90,-243)(613,-243)(613,79){7}
//: {8}(611,81)(607,81){9}
//: {10}(613,83)(613,91){11}
//: {12}(611,93)(607,93){13}
//: {14}(613,95)(613,104){15}
//: {16}(611,106)(607,106){17}
//: {18}(613,108)(613,116){19}
//: {20}(611,118)(607,118){21}
//: {22}(613,120)(613,128){23}
//: {24}(611,130)(607,130){25}
//: {26}(613,132)(-1:613,141){27}
//: {28}(611,143)(607,143){29}
//: {30}(613,145)(613,156)(607,156){31}
//: {32}(88,688)(70,688)(70,688)(61,688){33}
wire w23;    //: /sn:0 {0}(418,1685)(468,1685)(468,1647)(489,1647){1}
wire w298;    //: /sn:0 {0}(267,1205)(279,1205){1}
//: {2}(281,1203)(281,1175)(311,1175)(311,988){3}
//: {4}(313,986)(410,986)(410,986)(547,986){5}
//: {6}(311,984)(311,684)(990,684)(990,432)(778,432)(778,421){7}
//: {8}(780,419)(784,419){9}
//: {10}(776,419)(769,419)(769,411){11}
//: {12}(771,409)(774,409){13}
//: {14}(767,409)(760,409)(760,401){15}
//: {16}(762,399)(764,399){17}
//: {18}(758,399)(749,399)(749,390){19}
//: {20}(751,388)(755,388){21}
//: {22}(747,388)(741,388)(741,379){23}
//: {24}(743,377)(746,377){25}
//: {26}(739,377)(731,377)(731,369){27}
//: {28}(733,367)(735,367){29}
//: {30}(729,367)(722,367)(722,358){31}
//: {32}(724,356)(726,356){33}
//: {34}(720,356)(712,356)(712,347){35}
//: {36}(714,345)(716,345){37}
//: {38}(710,345)(703,345)(703,336){39}
//: {40}(705,334)(707,334){41}
//: {42}(701,334)(694,334)(694,325){43}
//: {44}(696,323)(697,323){45}
//: {46}(692,323)(686,323)(686,312)(688,312){47}
//: {48}(281,1207)(281,1256)(-500,1256)(-500,1340)(-490,1340){49}
wire w369;    //: /sn:0 {0}(-53,1370)(-60,1370){1}
wire w225;    //: /sn:0 {0}(535,1961)(530,1961){1}
wire w108;    //: /sn:0 {0}(547,1336)(451,1336)(451,1336)(396,1336){1}
//: {2}(394,1334)(394,609)(196,609)(196,-157)(562,-157)(562,-60){3}
//: {4}(560,-58)(559,-58)(559,-58)(558,-58){5}
//: {6}(562,-56)(562,-54)(563,-54)(563,-48){7}
//: {8}(561,-46)(560,-46){9}
//: {10}(563,-44)(563,-39)(565,-39)(565,-35){11}
//: {12}(563,-33)(560,-33)(560,-33)(562,-33){13}
//: {14}(565,-31)(565,-26)(568,-26)(568,-22){15}
//: {16}(566,-20)(565,-20)(565,-20)(565,-20){17}
//: {18}(568,-18)(568,-14)(571,-14)(571,-9){19}
//: {20}(569,-7)(568,-7){21}
//: {22}(571,-5)(571,-1)(573,-1)(573,3){23}
//: {24}(571,5)(571,5)(571,5)(570,5){25}
//: {26}(573,7)(573,12)(575,12)(575,16){27}
//: {28}(573,18)(572,18)(572,18)(572,18){29}
//: {30}(575,20)(575,24)(578,24)(578,29){31}
//: {32}(576,31)(575,31)(575,31)(575,31){33}
//: {34}(578,33)(578,37)(580,37)(580,41){35}
//: {36}(578,43)(577,43)(577,43)(577,43){37}
//: {38}(580,45)(580,50)(582,50)(582,54){39}
//: {40}(580,56)(579,56){41}
//: {42}(584,56)(587,56)(587,69)(582,69){43}
//: {44}(394,1338)(394,1614)(212,1614)(212,1641){45}
//: {46}(214,1643)(223,1643){47}
//: {48}(210,1643)(202,1643){49}
wire w300;    //: /sn:0 {0}(547,1056)(419,1056)(419,1056)(331,1056){1}
//: {2}(329,1054)(329,665)(589,665)(589,470){3}
//: {4}(591,468)(597,468)(597,468)(592,468){5}
//: {6}(589,466)(589,458){7}
//: {8}(591,456)(597,456)(597,456)(592,456){9}
//: {10}(589,454)(589,445){11}
//: {12}(591,443)(597,443)(597,443)(592,443){13}
//: {14}(589,441)(589,432){15}
//: {16}(591,430)(597,430)(597,430)(592,430){17}
//: {18}(589,428)(589,419)(589,419)(589,419){19}
//: {20}(591,417)(597,417)(597,417)(592,417){21}
//: {22}(589,415)(589,407){23}
//: {24}(591,405)(597,405)(597,405)(592,405){25}
//: {26}(589,403)(589,394){27}
//: {28}(591,392)(597,392)(597,392)(592,392){29}
//: {30}(589,390)(589,382){31}
//: {32}(591,380)(597,380)(597,380)(592,380){33}
//: {34}(589,378)(589,370){35}
//: {36}(591,368)(597,368)(597,368)(592,368){37}
//: {38}(589,366)(589,357){39}
//: {40}(591,355)(597,355)(597,355)(592,355){41}
//: {42}(589,353)(589,342)(592,342){43}
//: {44}(329,1058)(329,1290)(-47,1290)(-47,1345){45}
//: {46}(-45,1347)(-37,1347){47}
//: {48}(-49,1347)(-60,1347){49}
wire w223;    //: /sn:0 {0}(1056,1969)(1051,1969){1}
wire w125;    //: /sn:0 {0}(-62,824)(-69,824){1}
wire w8;    //: /sn:0 {0}(66,1904)(-900,1904)(-900,801)(-884,801){1}
wire w103;    //: /sn:0 {0}(547,866)(318,866)(318,866)(283,866){1}
//: {2}(281,864)(281,662)(147,662)(147,-197)(994,-197)(994,106)(865,106)(865,114)(855,114){3}
//: {4}(853,112)(853,111)(853,111)(853,110){5}
//: {6}(851,114)(849,114)(849,118)(844,118){7}
//: {8}(842,116)(842,115){9}
//: {10}(840,118)(835,118)(835,123)(831,123){11}
//: {12}(829,121)(829,118)(829,118)(829,120){13}
//: {14}(827,123)(822,123)(822,129)(818,129){15}
//: {16}(816,127)(816,126)(816,126)(816,126){17}
//: {18}(814,129)(810,129)(810,134)(806,134){19}
//: {20}(804,132)(804,131){21}
//: {22}(802,134)(798,134)(798,139)(794,139){23}
//: {24}(792,137)(792,137)(792,137)(792,136){25}
//: {26}(790,139)(785,139)(785,144)(781,144){27}
//: {28}(779,142)(779,141)(779,141)(779,141){29}
//: {30}(777,144)(773,144)(773,149)(769,149){31}
//: {32}(767,147)(767,146)(767,146)(767,146){33}
//: {34}(765,149)(761,149)(761,154)(757,154){35}
//: {36}(755,152)(755,151)(755,151)(755,151){37}
//: {38}(753,154)(748,154)(748,159)(744,159){39}
//: {40}(742,157)(742,156){41}
//: {42}(742,161)(742,164)(729,164)(729,161){43}
//: {44}(281,868)(281,881)(281,881)(281,1060){45}
//: {46}(279,1062)(267,1062){47}
//: {48}(281,1064)(281,1113)(-499,1113)(-499,1193)(-489,1193){49}
wire w202;    //: /sn:0 {0}(-363,1489)(-375,1489){1}
//: {2}(-377,1487)(-377,1415)(347,1415)(347,1128){3}
//: {4}(349,1126)(428,1126)(428,1126)(547,1126){5}
//: {6}(347,1124)(347,651)(297,651)(297,417)(403,417){7}
//: {8}(407,417)(409,417){9}
//: {10}(405,415)(405,406)(412,406){11}
//: {12}(416,406)(418,406)(418,406)(418,406){13}
//: {14}(414,404)(414,395)(420,395){15}
//: {16}(424,395)(427,395)(427,395)(427,395){17}
//: {18}(422,393)(422,384)(428,384){19}
//: {20}(432,384)(436,384)(436,384)(436,384){21}
//: {22}(430,382)(430,373)(438,373){23}
//: {24}(442,373)(445,373)(445,373)(445,373){25}
//: {26}(440,371)(440,362)(448,362){27}
//: {28}(452,362)(454,362)(454,362)(454,362){29}
//: {30}(1:450,360)(450,351)(457,351){31}
//: {32}(461,351)(463,351)(463,351)(463,351){33}
//: {34}(459,349)(459,340)(466,340){35}
//: {36}(470,340)(472,340)(472,340)(472,340){37}
//: {38}(468,338)(468,329)(472,329){39}
//: {40}(476,329)(480,329)(480,329)(481,329){41}
//: {42}(474,327)(474,318)(483,318){43}
//: {44}(487,318)(490,318)(490,318)(490,318){45}
//: {46}(485,316)(485,308)(499,308){47}
//: {48}(-379,1489)(-384,1489){49}
wire w314;    //: /sn:0 {0}(-295,1343)(-304,1343){1}
//: {2}(-306,1341)(-306,1274)(321,1274)(321,1018){3}
//: {4}(323,1016)(415,1016)(415,1016)(547,1016){5}
//: {6}(321,1014)(321,673)(688,673)(688,460){7}
//: {8}(690,458)(691,458)(691,458)(692,458){9}
//: {10}(688,456)(688,454)(684,454)(684,449){11}
//: {12}(686,447)(687,447){13}
//: {14}(684,445)(684,440)(679,440)(679,436){15}
//: {16}(681,434)(684,434)(684,434)(682,434){17}
//: {18}(679,432)(679,427)(673,427)(673,423){19}
//: {20}(675,421)(676,421)(676,421)(676,421){21}
//: {22}(673,419)(673,415)(668,415)(668,411){23}
//: {24}(670,409)(671,409){25}
//: {26}(668,407)(668,403)(663,403)(663,399){27}
//: {28}(665,397)(665,397)(665,397)(666,397){29}
//: {30}(663,395)(663,390)(658,390)(658,386){31}
//: {32}(660,384)(661,384)(661,384)(661,384){33}
//: {34}(658,382)(658,378)(653,378)(653,374){35}
//: {36}(655,372)(656,372)(656,372)(656,372){37}
//: {38}(653,370)(653,366)(648,366)(648,362){39}
//: {40}(650,360)(651,360)(651,360)(651,360){41}
//: {42}(648,358)(648,353)(643,353)(643,349){43}
//: {44}(645,347)(646,347){45}
//: {46}(641,347)(638,347)(638,334)(641,334){47}
//: {48}(-308,1343)(-321,1343){49}
wire w71;    //: /sn:0 {0}(224,1351)(221,1351){1}
//: {2}(219,1349)(219,1307)(337,1307)(337,1098){3}
//: {4}(339,1096)(423,1096)(423,1096)(547,1096){5}
//: {6}(337,1094)(337,657)(490,657)(490,459){7}
//: {8}(492,457)(492,457)(492,457)(492,457){9}
//: {10}(490,455)(490,451)(493,451)(493,447){11}
//: {12}(495,445)(496,445){13}
//: {14}(493,443)(493,438)(498,438)(498,435){15}
//: {16}(500,433)(505,433)(505,433)(501,433){17}
//: {18}(498,431)(498,426)(502,426)(502,422){19}
//: {20}(504,420)(511,420)(511,420)(507,420){21}
//: {22}(502,418)(502,409)(507,409)(507,410){23}
//: {24}(509,408)(516,408)(516,408)(512,408){25}
//: {26}(507,406)(507,402)(511,402)(511,397){27}
//: {28}(513,395)(520,395)(520,395)(516,395){29}
//: {30}(511,393)(511,388)(516,388)(516,385){31}
//: {32}(518,383)(525,383)(525,383)(521,383){33}
//: {34}(516,381)(516,377)(520,377)(520,373){35}
//: {36}(522,371)(529,371)(529,371)(525,371){37}
//: {38}(520,369)(520,365)(526,365)(526,361){39}
//: {40}(528,359)(535,359)(535,359)(531,359){41}
//: {42}(526,357)(526,352)(530,352)(530,349){43}
//: {44}(532,347)(539,347)(539,347)(535,347){45}
//: {46}(530,345)(530,334)(540,334){47}
//: {48}(217,1351)(203,1351){49}
wire w17;    //: /sn:0 {0}(-632,1060)(-642,1060)(-642,1888)(66,1888){1}
wire w297;    //: /sn:0 {0}(31,1348)(22,1348){1}
//: {2}(20,1346)(20,1294)(331,1294)(331,1068){3}
//: {4}(333,1066)(420,1066)(420,1066)(547,1066){5}
//: {6}(331,1064)(331,663)(561,663)(561,470){7}
//: {8}(563,468)(566,468){9}
//: {10}(561,466)(561,462)(563,462)(563,458){11}
//: {12}(565,456)(572,456)(572,456)(568,456){13}
//: {14}(563,454)(563,449)(564,449)(564,445){15}
//: {16}(566,443)(573,443)(573,443)(569,443){17}
//: {18}(564,441)(564,436)(566,436)(566,432){19}
//: {20}(568,430)(575,430)(575,430)(571,430){21}
//: {22}(566,428)(566,419)(567,419)(567,419){23}
//: {24}(569,417)(576,417)(576,417)(572,417){25}
//: {26}(567,415)(567,411)(568,411)(568,406){27}
//: {28}(570,404)(577,404)(577,404)(573,404){29}
//: {30}(568,402)(568,397)(569,397)(569,393){31}
//: {32}(571,391)(578,391)(578,391)(574,391){33}
//: {34}(569,389)(569,385)(570,385)(570,381){35}
//: {36}(572,379)(579,379)(579,379)(575,379){37}
//: {38}(570,377)(570,373)(571,373)(571,369){39}
//: {40}(573,367)(580,367)(580,367)(576,367){41}
//: {42}(571,365)(571,360)(573,360)(573,356){43}
//: {44}(575,354)(582,354)(582,354)(578,354){45}
//: {46}(573,352)(573,341)(579,341){47}
//: {48}(18,1348)(5,1348){49}
wire w84;    //: /sn:0 {0}(748,2233)(738,2233){1}
//: {2}(736,2231)(736,2175)(1360,2175)(1360,1276){3}
//: {4}(1360,1272)(1360,564)(211,564)(211,27)(359,27)(359,30){5}
//: {6}(1358,1274)(1197,1274){7}
//: {8}(734,2233)(724,2233){9}
wire w53;    //: /sn:0 {0}(615,1939)(606,1939){1}
//: {2}(604,1937)(604,1865)(1302,1865)(1302,1016){3}
//: {4}(1302,1012)(1302,625)(717,625)(717,461)(722,461){5}
//: {6}(1300,1014)(1197,1014){7}
//: {8}(602,1939)(594,1939){9}
wire w211;    //: /sn:0 {0}(97,1496)(86,1496){1}
//: {2}(84,1494)(84,1450)(361,1450)(361,1198){3}
//: {4}(363,1196)(435,1196)(435,1196)(547,1196){5}
//: {6}(361,1194)(361,641)(163,641)(163,216)(335,216){7}
//: {8}(339,216)(343,216)(343,215)(347,215){9}
//: {10}(349,217)(349,218){11}
//: {12}(351,215)(356,215)(356,214)(360,214){13}
//: {14}(362,216)(362,219)(362,219)(362,217){15}
//: {16}(364,214)(369,214)(369,213)(373,213){17}
//: {18}(375,215)(375,216)(375,216)(375,216){19}
//: {20}(377,213)(382,213)(382,212)(386,212){21}
//: {22}(388,214)(388,215){23}
//: {24}(390,212)(394,212)(394,211)(398,211){25}
//: {26}(400,213)(400,214)(400,214)(400,214){27}
//: {28}(402,211)(407,211)(407,210)(411,210){29}
//: {30}(413,212)(413,213)(413,213)(413,213){31}
//: {32}(415,210)(419,210)(419,209)(423,209){33}
//: {34}(425,211)(425,212)(425,212)(425,212){35}
//: {36}(427,209)(431,209)(431,208)(435,208){37}
//: {38}(437,210)(437,211)(437,211)(437,211){39}
//: {40}(439,208)(444,208)(444,207)(448,207){41}
//: {42}(450,209)(450,210){43}
//: {44}(452,207)(463,207)(463,209){45}
//: {46}(337,218)(337,219){47}
//: {48}(82,1496)(73,1496){49}
wire w2;    //: /sn:0 {0}(-653,1170)(-653,1040)(-632,1040){1}
wire w44;    //: /sn:0 {0}(792,1795)(801,1795){1}
//: {2}(805,1795)(814,1795){3}
//: {4}(803,1793)(803,1737)(1280,1737)(1280,926){5}
//: {6}(1280,922)(1280,649)(1033,649)(1033,248)(876,248)(876,237){7}
//: {8}(1278,924)(1197,924){9}
wire w113;    //: /sn:0 {0}(547,1026)(416,1026)(416,1026)(325,1026){1}
//: {2}(323,1024)(323,671)(662,671)(662,466){3}
//: {4}(664,464)(666,464){5}
//: {6}(662,462)(662,460)(660,460)(660,454){7}
//: {8}(662,452)(663,452){9}
//: {10}(660,450)(660,445)(656,445)(656,441){11}
//: {12}(658,439)(661,439)(661,439)(659,439){13}
//: {14}(656,437)(656,432)(652,432)(652,428){15}
//: {16}(654,426)(655,426)(655,426)(655,426){17}
//: {18}(652,424)(652,420)(648,420)(648,415){19}
//: {20}(650,413)(651,413){21}
//: {22}(648,411)(648,407)(645,407)(645,403){23}
//: {24}(647,401)(647,401)(647,401)(648,401){25}
//: {26}(645,399)(645,394)(641,394)(641,391){27}
//: {28}(643,389)(644,389)(644,389)(644,389){29}
//: {30}(641,387)(641,383)(637,383)(637,378){31}
//: {32}(639,376)(640,376)(640,376)(640,376){33}
//: {34}(637,374)(637,370)(634,370)(634,366){35}
//: {36}(636,364)(637,364)(637,364)(637,364){37}
//: {38}(634,362)(634,357)(630,357)(630,353){39}
//: {40}(632,351)(633,351){41}
//: {42}(628,351)(625,351)(625,338)(629,338){43}
//: {44}(323,1028)(323,1278)(-241,1278)(-241,1342){45}
//: {46}(-239,1344)(-229,1344){47}
//: {48}(-243,1344)(-253,1344){49}
wire w345;    //: /sn:0 {0}(-441,1074)(-447,1074){1}
wire fdbk60;    //: /sn:0 {0}(-616,1073)(-616,1088){1}
//: {2}(-618,1090)(-837,1090)(-837,895){3}
//: {4}(-837,891)(-837,881)(-837,881)(-837,871){5}
//: {6}(-839,893)(-868,893)(-868,814){7}
//: {8}(-616,1092)(-616,1139)(-616,1139)(-616,1149){9}
//: {10}(-614,1151)(-588,1151)(-588,1131){11}
//: {12}(-616,1153)(-616,1755)(234,1755){13}
//: {14}(238,1755)(316,1755)(316,1780)(304,1780){15}
//: {16}(236,1757)(236,1866)(197,1866){17}
wire w83;    //: /sn:0 {0}(682,2232)(672,2232){1}
//: {2}(670,2230)(670,2170)(1358,2170)(1358,1266){3}
//: {4}(1358,1262)(1358,566)(209,566)(209,58)(346,58)(346,67){5}
//: {6}(1356,1264)(1197,1264){7}
//: {8}(668,2232)(656,2232){9}
wire w77;    //: /sn:0 {0}(1181,2095)(1189,2095){1}
//: {2}(1193,2095)(1202,2095){3}
//: {4}(1191,2093)(1191,2057)(1347,2057)(1347,1226){5}
//: {6}(1347,1222)(1347,579)(236,579)(236,161)(322,161)(322,168){7}
//: {8}(1345,1224)(1197,1224){9}
wire w367;    //: /sn:0 {0}(-314,1513)(-321,1513){1}
wire w224;    //: /sn:0 {0}(-296,1635)(-306,1635){1}
//: {2}(-308,1633)(-308,1573)(378,1573)(378,1258){3}
//: {4}(380,1256)(443,1256)(443,1256)(547,1256){5}
//: {6}(378,1254)(378,625)(180,625)(180,63)(358,63){7}
//: {8}(362,63)(372,63)(372,67){9}
//: {10}(374,69)(384,69)(384,72){11}
//: {12}(386,74)(396,74)(396,78){13}
//: {14}(396,82)(396,91){15}
//: {16}(398,80)(408,80)(408,84){17}
//: {18}(408,88)(408,97){19}
//: {20}(410,86)(420,86)(420,92){21}
//: {22}(420,96)(420,103){23}
//: {24}(422,94)(1:432,94)(432,100){25}
//: {26}(432,104)(432,109){27}
//: {28}(434,102)(444,102)(444,102){29}
//: {30}(444,106)(444,114){31}
//: {32}(446,104)(456,104)(456,108){33}
//: {34}(456,112)(456,120){35}
//: {36}(458,110)(468,110)(468,113){37}
//: {38}(468,117)(468,126){39}
//: {40}(470,115)(480,115)(480,132){41}
//: {42}(384,76)(384,85){43}
//: {44}(372,71)(372,79){45}
//: {46}(360,65)(360,73){47}
//: {48}(-310,1635)(-322,1635){49}
wire w274;    //: /sn:0 {0}(161,1497)(154,1497){1}
//: {2}(152,1495)(152,1456)(363,1456)(363,1208){3}
//: {4}(365,1206)(436,1206)(436,1206)(547,1206){5}
//: {6}(363,1204)(363,639)(165,639)(165,192)(335,192){7}
//: {8}(339,192)(347,192){9}
//: {10}(349,194)(349,200)(349,200)(349,195){11}
//: {12}(351,192)(360,192){13}
//: {14}(362,194)(362,200)(362,200)(362,195){15}
//: {16}(364,192)(373,192){17}
//: {18}(375,194)(375,200)(375,200)(375,195){19}
//: {20}(377,192)(386,192)(386,192)(386,192){21}
//: {22}(388,194)(388,200)(388,200)(388,195){23}
//: {24}(390,192)(398,192){25}
//: {26}(400,194)(400,200)(400,200)(400,195){27}
//: {28}(402,192)(411,192){29}
//: {30}(413,194)(413,200)(413,200)(413,195){31}
//: {32}(415,192)(423,192){33}
//: {34}(425,194)(425,200)(425,200)(425,195){35}
//: {36}(427,192)(435,192){37}
//: {38}(439,192)(448,192){39}
//: {40}(450,194)(450,200)(450,200)(450,195){41}
//: {42}(452,192)(463,192)(463,195){43}
//: {44}(437,194)(437,200)(437,200)(437,195){45}
//: {46}(337,194)(337,200)(337,200)(337,195){47}
//: {48}(150,1497)(139,1497){49}
wire w366;    //: /sn:0 {0}(-376,1218)(-383,1218){1}
wire w362;    //: /sn:0 {0}(79,1225)(74,1225){1}
wire w351;    //: /sn:0 {0}(145,1083)(140,1083){1}
wire w315;    //: /sn:0 {0}(-52,1223)(-59,1223){1}
wire w262;    //: /sn:0 {0}(861,2258)(854,2258){1}
wire w10;    //: /sn:0 {0}(814,1652)(807,1652){1}
//: {2}(805,1650)(805,1524)(1252,1524)(1252,806){3}
//: {4}(1252,802)(1252,681)(1013,681)(1013,-181)(758,-181)(758,-61)(714,-61){5}
//: {6}(1250,804)(1197,804){7}
//: {8}(803,1652)(792,1652){9}
wire w275;    //: /sn:0 {0}(534,2253)(529,2253){1}
wire w273;    //: /sn:0 {0}(1055,2261)(1050,2261){1}
wire w95;    //: /sn:0 {0}(982,2237)(996,2237){1}
//: {2}(1000,2237)(1008,2237){3}
//: {4}(998,2235)(998,2195)(1368,2195)(1368,1316){5}
//: {6}(1368,1312)(1368,556)(219,556)(219,-170)(485,-170)(485,-54)(479,-54){7}
//: {8}(1366,1314)(1197,1314){9}
wire w52;    //: /sn:0 {0}(488,1937)(478,1937)(478,1853)(1259,1853)(1259,1804){1}
//: {2}(1259,1800)(1259,1763)(1294,1763)(1294,996){3}
//: {4}(1294,992)(1294,629)(788,629)(788,431)(794,431){5}
//: {6}(1292,994)(1197,994){7}
//: {8}(1257,1802)(1245,1802){9}
wire w178;    //: /sn:0 {0}(1123,1823)(1118,1823){1}
wire w50;    //: /sn:0 {0}(1118,1800)(1128,1800){1}
//: {2}(1132,1800)(1140,1800){3}
//: {4}(1130,1798)(1130,1756)(1290,1756)(1290,976){5}
//: {6}(1290,972)(1290,639)(1043,639)(1043,380)(843,380)(843,377){7}
//: {8}(1288,974)(1197,974){9}
wire w330;    //: /sn:0 {0}(-425,1194)(-433,1194){1}
//: {2}(-435,1192)(-435,1129)(289,1129)(289,878){3}
//: {4}(291,876)(399,876)(399,876)(547,876){5}
//: {6}(289,874)(289,655)(149,655)(149,-195)(992,-195)(992,150)(859,150)(859,142){7}
//: {8}(859,138)(859,137)(859,137)(859,136){9}
//: {10}(857,140)(855,140)(855,142)(849,142){11}
//: {12}(847,140)(847,139){13}
//: {14}(845,142)(840,142)(840,146)(836,146){15}
//: {16}(834,144)(834,141)(834,141)(834,143){17}
//: {18}(832,146)(827,146)(827,150)(823,150){19}
//: {20}(821,148)(821,147)(821,147)(821,147){21}
//: {22}(819,150)(815,150)(815,154)(810,154){23}
//: {24}(808,152)(808,151){25}
//: {26}(806,154)(802,154)(802,157)(798,157){27}
//: {28}(796,155)(796,155)(796,155)(796,154){29}
//: {30}(794,157)(789,157)(789,161)(786,161){31}
//: {32}(784,159)(784,158)(784,158)(784,158){33}
//: {34}(782,161)(778,161)(778,165)(773,165){35}
//: {36}(771,163)(771,162)(771,162)(771,162){37}
//: {38}(769,165)(765,165)(765,168)(761,168){39}
//: {40}(759,166)(759,165)(759,165)(759,165){41}
//: {42}(757,168)(752,168)(752,172)(748,172){43}
//: {44}(746,170)(746,169){45}
//: {46}(746,174)(746,177)(733,177)(733,173){47}
//: {48}(-437,1194)(-447,1194){49}
wire w6;    //: /sn:0 {0}(684,1650)(669,1650){1}
//: {2}(667,1648)(667,1516)(1248,1516)(1248,786){3}
//: {4}(1248,782)(1248,685)(1017,685)(1017,-185)(688,-185)(688,-72)(661,-72){5}
//: {6}(1246,784)(1197,784){7}
//: {8}(665,1650)(658,1650){9}
wire w93;    //: /sn:0 {0}(790,2234)(800,2234){1}
//: {2}(804,2234)(812,2234){3}
//: {4}(802,2232)(802,2180)(1362,2180)(1362,1286){5}
//: {6}(1362,1282)(1362,562)(213,562)(213,-164)(375,-164)(375,0){7}
//: {8}(1360,1284)(1197,1284){9}
wire w7;    //: /sn:0 {0}(66,1872)(56,1872){1}
//: {2}(54,1870)(54,1847)(218,1847)(218,1874)(291,1874)(291,1856){3}
//: {4}(291,1852)(291,1796){5}
//: {6}(289,1854)(268,1854)(268,1823){7}
//: {8}(52,1872)(-656,1872)(-656,1191){9}
wire w61;    //: /sn:0 {0}(-603,1050)(-564,1050)(-564,1050)(-552,1050){1}
//: {2}(-548,1050)(-517,1050)(-517,1050)(-489,1050){3}
//: {4}(-550,1048)(-550,1038)(-550,1038)(-550,992){5}
wire w99;    //: /sn:0 {0}(665,1673)(658,1673){1}
wire w153;    //: /sn:0 {0}(-101,1056)(-111,1056){1}
//: {2}(-113,1054)(-113,932)(269,932)(269,808){3}
//: {4}(271,806)(299,806)(299,806)(547,806){5}
//: {6}(269,804)(269,674)(135,674)(135,-209)(740,-209)(740,-39){7}
//: {8}(738,-37)(730,-37){9}
//: {10}(740,-35)(740,-25)(736,-25){11}
//: {12}(732,-25)(724,-25){13}
//: {14}(734,-23)(734,-13)(731,-13){15}
//: {16}(727,-13)(718,-13){17}
//: {18}(729,-11)(729,-1)(725,-1){19}
//: {20}(721,-1)(712,-1){21}
//: {22}(723,1)(723,11)(719,11){23}
//: {24}(715,11)(706,11){25}
//: {26}(717,13)(717,23)(711,23){27}
//: {28}(707,23)(700,23){29}
//: {30}(709,25)(1:709,35)(703,35){31}
//: {32}(699,35)(694,35){33}
//: {34}(701,37)(701,47)(701,47){35}
//: {36}(697,47)(689,47){37}
//: {38}(699,49)(699,59)(695,59){39}
//: {40}(691,59)(683,59){41}
//: {42}(693,61)(693,71)(690,71){43}
//: {44}(686,71)(677,71){45}
//: {46}(688,73)(688,83)(671,83){47}
//: {48}(-115,1056)(-122,1056){49}
wire w135;    //: /sn:0 {0}(1252,2264)(1243,2264){1}
wire w352;    //: /sn:0 {0}(349,147)(349,151)(349,151)(349,145){1}
//: {2}(347,143)(343,143)(343,140)(339,140){3}
//: {4}(335,140)(169,140)(169,635)(367,635)(367,1224){5}
//: {6}(369,1226)(438,1226)(438,1226)(547,1226){7}
//: {8}(367,1228)(367,1468)(280,1468)(280,1497){9}
//: {10}(278,1499)(266,1499){11}
//: {12}(280,1501)(280,1551)(-501,1551)(-501,1632)(-491,1632){13}
//: {14}(337,142)(337,148)(337,148)(337,144){15}
//: {16}(351,143)(356,143)(356,145)(360,145){17}
//: {18}(362,147)(362,153)(362,153)(362,149){19}
//: {20}(364,145)(369,145)(369,147)(373,147){21}
//: {22}(375,149)(375,156)(375,156)(375,152){23}
//: {24}(377,147)(386,147)(386,150)(386,150){25}
//: {26}(388,152)(388,159)(388,159)(388,155){27}
//: {28}(390,150)(394,150)(394,152)(399,152){29}
//: {30}(401,154)(401,161)(401,161)(401,157){31}
//: {32}(403,152)(408,152)(408,154)(412,154){33}
//: {34}(414,156)(414,163)(414,163)(414,159){35}
//: {36}(416,154)(420,154)(420,156)(424,156){37}
//: {38}(426,158)(426,165)(426,165)(426,161){39}
//: {40}(428,156)(432,156)(432,159)(436,159){41}
//: {42}(438,161)(438,168)(438,168)(438,164){43}
//: {44}(440,159)(445,159)(445,162)(449,162){45}
//: {46}(451,164)(451,171)(451,171)(451,167){47}
//: {48}(453,162)(464,162)(464,169){49}
wire w380;    //: /sn:0 {0}(273,1522)(266,1522){1}
wire w288;    //: /sn:0 {0}(211,1227)(204,1227){1}
wire w51;    //: /sn:0 {0}(1182,1801)(1192,1801){1}
//: {2}(1196,1801)(1203,1801){3}
//: {4}(1194,1799)(1194,1759)(1292,1759)(1292,986){5}
//: {6}(1292,982)(1292,637)(1045,637)(1045,415)(826,415)(826,408){7}
//: {8}(1290,984)(1197,984){9}
wire w207;    //: /sn:0 {0}(547,1166)(432,1166)(432,1166)(357,1166){1}
//: {2}(355,1164)(355,647)(157,647)(157,292)(345,292){3}
//: {4}(349,292)(351,292)(351,288)(356,288){5}
//: {6}(358,290)(358,291){7}
//: {8}(360,288)(365,288)(365,283)(369,283){9}
//: {10}(371,285)(371,288)(371,288)(371,286){11}
//: {12}(373,283)(378,283)(378,277)(382,277){13}
//: {14}(384,279)(384,280)(384,280)(384,280){15}
//: {16}(386,277)(390,277)(390,272)(394,272){17}
//: {18}(396,274)(396,275){19}
//: {20}(398,272)(402,272)(402,267)(406,267){21}
//: {22}(408,269)(408,269)(408,269)(408,270){23}
//: {24}(410,267)(415,267)(415,262)(419,262){25}
//: {26}(421,264)(421,265)(421,265)(421,265){27}
//: {28}(423,262)(427,262)(427,257)(431,257){29}
//: {30}(433,259)(433,260)(433,260)(433,260){31}
//: {32}(435,257)(439,257)(439,252)(443,252){33}
//: {34}(445,254)(445,255)(445,255)(445,255){35}
//: {36}(447,252)(452,252)(452,247)(456,247){37}
//: {38}(458,249)(458,250){39}
//: {40}(458,245)(458,242)(471,242)(471,245){41}
//: {42}(347,294)(347,295)(347,295)(347,296){43}
//: {44}(355,1168)(355,1435)(-117,1435)(-117,1491){45}
//: {46}(-115,1493)(-102,1493){47}
//: {48}(-119,1493)(-123,1493){49}
wire w239;    //: /sn:0 {0}(730,2111)(725,2111){1}
wire w106;    //: /sn:0 {0}(1252,1682)(1245,1682){1}
wire w304;    //: /sn:0 {0}(547,1086)(422,1086)(422,1086)(337,1086){1}
//: {2}(335,1084)(335,659)(513,659)(513,468){3}
//: {4}(515,466)(516,466){5}
//: {6}(513,464)(513,460)(517,460)(517,456){7}
//: {8}(519,454)(524,454)(524,454)(520,454){9}
//: {10}(517,452)(517,447)(520,447)(520,443){11}
//: {12}(522,441)(527,441)(527,441)(523,441){13}
//: {14}(520,439)(520,434)(523,434)(523,430){15}
//: {16}(525,428)(532,428)(532,428)(528,428){17}
//: {18}(523,426)(523,417)(527,417)(527,417){19}
//: {20}(529,415)(536,415)(536,415)(532,415){21}
//: {22}(527,413)(527,409)(530,409)(530,404){23}
//: {24}(532,402)(539,402)(539,402)(535,402){25}
//: {26}(530,400)(530,395)(533,395)(533,391){27}
//: {28}(535,389)(542,389)(542,389)(538,389){29}
//: {30}(533,387)(533,383)(536,383)(536,379){31}
//: {32}(538,377)(545,377)(545,377)(541,377){33}
//: {34}(536,375)(536,371)(541,371)(541,367){35}
//: {36}(543,365)(550,365)(550,365)(546,365){37}
//: {38}(541,363)(541,358)(545,358)(545,354){39}
//: {40}(547,352)(554,352)(554,352)(550,352){41}
//: {42}(545,350)(545,339)(553,339){43}
//: {44}(335,1088)(335,1302)(153,1302)(153,1348){45}
//: {46}(155,1350)(161,1350){47}
//: {48}(151,1350)(139,1350){49}
wire w373;    //: /sn:0 {0}(-443,1511)(-448,1511){1}
wire w349;    //: /sn:0 {0}(144,1520)(139,1520){1}
wire w69;    //: /sn:0 {0}(643,481)(631,481)(631,619)(1308,619)(1308,1042){1}
//: {2}(1306,1044)(1197,1044){3}
//: {4}(1308,1046)(1308,1878)(800,1878)(800,1940){5}
//: {6}(802,1942)(813,1942){7}
//: {8}(798,1942)(791,1942){9}
wire w357;    //: /sn:0 {0}(-164,1055)(-171,1055){1}
//: {2}(-173,1053)(-173,929)(267,929)(267,798){3}
//: {4}(269,796)(296,796)(296,796)(547,796){5}
//: {6}(267,794)(267,676)(133,676)(133,-211)(499,-211)(709,-211)(709,-49){7}
//: {8}(707,-47)(707,-47)(707,-47)(707,-47){9}
//: {10}(709,-45)(709,-41)(706,-41)(706,-37){11}
//: {12}(704,-35)(703,-35){13}
//: {14}(706,-33)(706,-28)(701,-28)(701,-25){15}
//: {16}(699,-23)(694,-23)(694,-23)(698,-23){17}
//: {18}(701,-21)(701,-16)(697,-16)(697,-12){19}
//: {20}(695,-10)(688,-10)(688,-10)(692,-10){21}
//: {22}(697,-8)(697,1)(692,1)(692,0){23}
//: {24}(690,2)(683,2)(683,2)(687,2){25}
//: {26}(692,4)(692,8)(688,8)(688,13){27}
//: {28}(686,15)(679,15)(679,15)(683,15){29}
//: {30}(688,17)(688,22)(683,22)(683,25){31}
//: {32}(681,27)(674,27)(674,27)(678,27){33}
//: {34}(683,29)(683,33)(679,33)(679,37){35}
//: {36}(677,39)(670,39)(670,39)(674,39){37}
//: {38}(679,41)(679,45)(673,45)(673,49){39}
//: {40}(671,51)(664,51)(664,51)(668,51){41}
//: {42}(673,53)(673,58)(669,58)(669,61){43}
//: {44}(667,63)(660,63)(660,63)(664,63){45}
//: {46}(669,65)(669,76)(659,76){47}
//: {48}(-175,1055)(-186,1055){49}
wire w177;    //: /sn:0 {0}(32,1201)(22,1201){1}
//: {2}(20,1199)(20,1158)(303,1158)(303,948){3}
//: {4}(305,946)(406,946)(406,946)(547,946){5}
//: {6}(303,944)(303,692)(982,692)(982,319)(851,319)(851,315){7}
//: {8}(851,311)(851,311)(851,311)(851,311){9}
//: {10}(849,313)(845,313)(845,310)(841,310){11}
//: {12}(839,308)(839,307){13}
//: {14}(837,310)(832,310)(832,305)(829,305){15}
//: {16}(827,303)(827,298)(827,298)(827,302){17}
//: {18}(825,305)(820,305)(820,301)(816,301){19}
//: {20}(814,299)(814,292)(814,292)(814,296){21}
//: {22}(812,301)(803,301)(803,296)(804,296){23}
//: {24}(802,294)(802,287)(802,287)(802,291){25}
//: {26}(800,296)(796,296)(796,292)(791,292){27}
//: {28}(789,290)(789,283)(789,283)(789,287){29}
//: {30}(787,292)(782,292)(782,287)(779,287){31}
//: {32}(777,285)(777,278)(777,278)(777,282){33}
//: {34}(775,287)(771,287)(771,283)(767,283){35}
//: {36}(765,281)(765,274)(765,274)(765,278){37}
//: {38}(763,283)(759,283)(759,277)(755,277){39}
//: {40}(753,275)(753,268)(753,268)(753,272){41}
//: {42}(751,277)(746,277)(746,273)(743,273){43}
//: {44}(741,271)(741,264)(741,264)(741,268){45}
//: {46}(739,273)(728,273)(728,263){47}
//: {48}(18,1201)(6,1201){49}
wire w66;    //: /sn:0 {0}(530,2085)(539,2085){1}
//: {2}(543,2085)(552,2085){3}
//: {4}(541,2083)(541,2003)(1327,2003)(1327,1126){5}
//: {6}(1327,1122)(1327,599)(256,599)(256,460)(421,460)(421,445)(429,445){7}
//: {8}(1325,1124)(1197,1124){9}
wire w290;    //: /sn:0 {0}(-364,1634)(-374,1634){1}
//: {2}(-376,1632)(-376,1567)(376,1567)(376,1248){3}
//: {4}(378,1246)(442,1246)(442,1246)(547,1246){5}
//: {6}(376,1244)(376,627)(178,627)(178,93)(346,93){7}
//: {8}(348,95)(348,95)(348,95)(348,95){9}
//: {10}(350,93)(354,93)(354,96)(358,96){11}
//: {12}(360,98)(360,99){13}
//: {14}(362,96)(367,96)(367,101)(370,101){15}
//: {16}(374,101)(379,101)(379,105)(383,105){17}
//: {18}(387,105)(396,105)(396,110)(395,110){19}
//: {20}(397,112)(397,119)(397,119)(397,115){21}
//: {22}(399,110)(403,110)(403,114)(408,114){23}
//: {24}(410,116)(410,123)(410,123)(410,119){25}
//: {26}(412,114)(417,114)(417,119)(420,119){27}
//: {28}(422,121)(422,128)(422,128)(422,124){29}
//: {30}(424,119)(428,119)(428,123)(432,123){31}
//: {32}(434,125)(434,132)(434,132)(434,128){33}
//: {34}(436,123)(440,123)(440,129)(444,129){35}
//: {36}(446,131)(446,138)(446,138)(446,134){37}
//: {38}(448,129)(453,129)(453,133)(456,133){39}
//: {40}(458,135)(458,142)(458,142)(458,138){41}
//: {42}(460,133)(471,133)(471,143){43}
//: {44}(385,107)(385,110){45}
//: {46}(372,103)(372,108)(372,108)(372,104){47}
//: {48}(-378,1634)(-385,1634){49}
wire [11:0] w37;    //: /sn:0 {0}(#:-94,584)(-100,584)(-100,633)(#:55,633){1}
wire w34;    //: /sn:0 {0}(225,1228)(216,1228)(216,1251)(152,1251){1}
//: {2}(150,1249)(150,1227)(162,1227){3}
//: {4}(148,1251)(136,1251)(136,1251)(90,1251){5}
//: {6}(88,1249)(88,1226)(98,1226){7}
//: {8}(86,1251)(55,1251)(55,1251)(23,1251){9}
//: {10}(21,1249)(21,1225)(32,1225){11}
//: {12}(19,1251)(-37,1251)(-37,1251)(-44,1251){13}
//: {14}(-46,1249)(-46,1224)(-36,1224){15}
//: {16}(-48,1251)(-59,1251)(-59,1251)(-109,1251){17}
//: {18}(-111,1249)(-111,1223)(-101,1223){19}
//: {20}(-113,1251)(-174,1251){21}
//: {22}(-176,1249)(-176,1222)(-164,1222){23}
//: {24}(-178,1251)(-190,1251)(-190,1251)(-236,1251){25}
//: {26}(-238,1249)(-238,1221)(-228,1221){27}
//: {28}(-240,1251)(-271,1251)(-271,1251)(-303,1251){29}
//: {30}(-305,1249)(-305,1220)(-294,1220){31}
//: {32}(-307,1251)(-363,1251)(-363,1251)(-370,1251){33}
//: {34}(-372,1249)(-372,1219)(-362,1219){35}
//: {36}(-374,1251)(-435,1251){37}
//: {38}(-437,1249)(-437,1218)(-425,1218){39}
//: {40}(-439,1251)(-451,1251)(-451,1251)(-497,1251){41}
//: {42}(-499,1249)(-499,1217)(-489,1217){43}
//: {44}(-501,1251)(-530,1251){45}
//: {46}(-532,1249)(-532,1110){47}
//: {48}(-530,1108)(-501,1108){49}
//: {50}(-497,1108)(-451,1108)(-451,1108)(-439,1108){51}
//: {52}(-435,1108)(-374,1108){53}
//: {54}(-370,1108)(-363,1108)(-363,1108)(-307,1108){55}
//: {56}(-303,1108)(-271,1108)(-271,1108)(-240,1108){57}
//: {58}(-236,1108)(-190,1108)(-190,1108)(-178,1108){59}
//: {60}(-174,1108)(-113,1108){61}
//: {62}(-109,1108)(-59,1108)(-59,1108)(-48,1108){63}
//: {64}(-44,1108)(-37,1108)(-37,1108)(19,1108){65}
//: {66}(23,1108)(55,1108)(55,1108)(86,1108){67}
//: {68}(90,1108)(136,1108)(136,1108)(148,1108){69}
//: {70}(152,1108)(182,1108)(182,1108)(216,1108)(216,1085)(225,1085){71}
//: {72}(150,1106)(150,1084)(162,1084){73}
//: {74}(88,1106)(88,1083)(98,1083){75}
//: {76}(21,1106)(21,1082)(32,1082){77}
//: {78}(-46,1106)(-46,1081)(-36,1081){79}
//: {80}(-111,1106)(-111,1080)(-101,1080){81}
//: {82}(-176,1106)(-176,1079)(-164,1079){83}
//: {84}(-238,1106)(-238,1078)(-228,1078){85}
//: {86}(-305,1106)(-305,1077)(-294,1077){87}
//: {88}(-372,1106)(-372,1076)(-362,1076){89}
//: {90}(-437,1106)(-437,1075)(-425,1075){91}
//: {92}(-499,1106)(-499,1074)(-489,1074){93}
//: {94}(-532,1106)(-532,940)(-517,940)(-517,925)(-527,925){95}
//: {96}(-532,1253)(-532,1396){97}
//: {98}(-530,1398)(-502,1398){99}
//: {100}(-498,1398)(-452,1398)(-452,1398)(-440,1398){101}
//: {102}(-436,1398)(-375,1398){103}
//: {104}(-371,1398)(-364,1398)(-364,1398)(-308,1398){105}
//: {106}(-304,1398)(-272,1398)(-272,1398)(-241,1398){107}
//: {108}(-237,1398)(-191,1398)(-191,1398)(-179,1398){109}
//: {110}(-175,1398)(-114,1398){111}
//: {112}(-110,1398)(-60,1398)(-60,1398)(-49,1398){113}
//: {114}(-45,1398)(-38,1398)(-38,1398)(18,1398){115}
//: {116}(22,1398)(54,1398)(54,1398)(85,1398){117}
//: {118}(89,1398)(135,1398)(135,1398)(147,1398){119}
//: {120}(151,1398)(181,1398)(181,1398)(215,1398)(215,1375)(224,1375){121}
//: {122}(149,1396)(149,1374)(161,1374){123}
//: {124}(87,1396)(87,1373)(97,1373){125}
//: {126}(20,1396)(20,1372)(31,1372){127}
//: {128}(-47,1396)(-47,1371)(-37,1371){129}
//: {130}(-112,1396)(-112,1370)(-102,1370){131}
//: {132}(-177,1396)(-177,1369)(-165,1369){133}
//: {134}(-239,1396)(-239,1368)(-229,1368){135}
//: {136}(-306,1396)(-306,1367)(-295,1367){137}
//: {138}(-373,1396)(-373,1366)(-363,1366){139}
//: {140}(-438,1396)(-438,1365)(-426,1365){141}
//: {142}(-500,1396)(-500,1364)(-490,1364){143}
//: {144}(-532,1400)(-532,1543){145}
//: {146}(-530,1545)(-502,1545){147}
//: {148}(-498,1545)(-452,1545)(-452,1545)(-440,1545){149}
//: {150}(-436,1545)(-375,1545){151}
//: {152}(-371,1545)(-364,1545)(-364,1545)(-308,1545){153}
//: {154}(-304,1545)(-272,1545)(-272,1545)(-241,1545){155}
//: {156}(-237,1545)(-191,1545)(-191,1545)(-179,1545){157}
//: {158}(-175,1545)(-114,1545){159}
//: {160}(-110,1545)(-60,1545)(-60,1545)(-49,1545){161}
//: {162}(-45,1545)(-38,1545)(-38,1545)(18,1545){163}
//: {164}(22,1545)(54,1545)(54,1545)(85,1545){165}
//: {166}(89,1545)(135,1545)(135,1545)(147,1545){167}
//: {168}(151,1545)(181,1545)(181,1545)(213,1545){169}
//: {170}(217,1545)(288,1545){171}
//: {172}(215,1543)(215,1522)(224,1522){173}
//: {174}(149,1543)(149,1521)(161,1521){175}
//: {176}(87,1543)(87,1520)(97,1520){177}
//: {178}(20,1543)(20,1519)(31,1519){179}
//: {180}(-47,1543)(-47,1518)(-37,1518){181}
//: {182}(-112,1543)(-112,1517)(-102,1517){183}
//: {184}(-177,1543)(-177,1516)(-165,1516){185}
//: {186}(-239,1543)(-239,1515)(-229,1515){187}
//: {188}(-306,1543)(-306,1514)(-295,1514){189}
//: {190}(-373,1543)(-373,1513)(-363,1513){191}
//: {192}(-438,1543)(-438,1512)(-426,1512){193}
//: {194}(-500,1543)(-500,1511)(-490,1511){195}
//: {196}(-532,1547)(-532,1690)(-503,1690){197}
//: {198}(-499,1690)(-453,1690)(-453,1690)(-441,1690){199}
//: {200}(-437,1690)(-376,1690){201}
//: {202}(-372,1690)(-365,1690)(-365,1690)(-309,1690){203}
//: {204}(-305,1690)(-273,1690)(-273,1690)(-242,1690){205}
//: {206}(-238,1690)(-192,1690)(-192,1690)(-180,1690){207}
//: {208}(-176,1690)(-115,1690){209}
//: {210}(-111,1690)(-61,1690)(-61,1690)(-50,1690){211}
//: {212}(-46,1690)(-39,1690)(-39,1690)(17,1690){213}
//: {214}(21,1690)(53,1690)(53,1690)(84,1690){215}
//: {216}(88,1690)(134,1690)(134,1690)(146,1690){217}
//: {218}(150,1690)(214,1690)(214,1667)(223,1667){219}
//: {220}(148,1688)(148,1666)(160,1666){221}
//: {222}(86,1688)(86,1665)(96,1665){223}
//: {224}(19,1688)(19,1664)(30,1664){225}
//: {226}(-48,1688)(-48,1663)(-38,1663){227}
//: {228}(-113,1688)(-113,1662)(-103,1662){229}
//: {230}(-178,1688)(-178,1661)(-166,1661){231}
//: {232}(-240,1688)(-240,1660)(-230,1660){233}
//: {234}(-307,1688)(-307,1659)(-296,1659){235}
//: {236}(-374,1688)(-374,1658)(-364,1658){237}
//: {238}(-439,1688)(-439,1657)(-427,1657){239}
//: {240}(-501,1688)(-501,1656)(-491,1656){241}
wire w299;    //: /sn:0 {0}(274,1228)(267,1228){1}
wire w356;    //: /sn:0 {0}(-37,1494)(-47,1494){1}
//: {2}(-49,1492)(-49,1440)(357,1440)(357,1178){3}
//: {4}(359,1176)(433,1176)(433,1176)(547,1176){5}
//: {6}(357,1174)(357,645)(159,645)(159,266)(339,266){7}
//: {8}(343,266)(345,266)(345,264)(351,264){9}
//: {10}(353,266)(353,267){11}
//: {12}(355,264)(360,264)(360,260)(364,260){13}
//: {14}(366,262)(366,265)(366,265)(366,263){15}
//: {16}(368,260)(373,260)(373,256)(377,256){17}
//: {18}(379,258)(379,259)(379,259)(379,259){19}
//: {20}(381,256)(385,256)(385,252)(390,252){21}
//: {22}(392,254)(392,255){23}
//: {24}(394,252)(398,252)(398,249)(402,249){25}
//: {26}(404,251)(404,251)(404,251)(404,252){27}
//: {28}(406,249)(411,249)(411,245)(414,245){29}
//: {30}(416,247)(416,248)(416,248)(416,248){31}
//: {32}(418,245)(422,245)(422,241)(427,241){33}
//: {34}(429,243)(429,244)(429,244)(429,244){35}
//: {36}(431,241)(435,241)(435,238)(439,238){37}
//: {38}(441,240)(441,241)(441,241)(441,241){39}
//: {40}(443,238)(448,238)(448,234)(452,234){41}
//: {42}(454,236)(454,237){43}
//: {44}(454,232)(454,229)(467,229)(467,233){45}
//: {46}(341,268)(341,269)(341,269)(341,270){47}
//: {48}(-51,1494)(-60,1494){49}
wire w87;    //: /sn:0 {0}(547,816)(305,816)(305,816)(273,816){1}
//: {2}(271,814)(271,672)(137,672)(137,-207)(777,-207)(777,-38)(769,-38)(769,-28){3}
//: {4}(767,-26)(764,-26){5}
//: {6}(769,-24)(769,-14)(764,-14){7}
//: {8}(760,-14)(757,-14){9}
//: {10}(762,-12)(762,-2)(757,-2){11}
//: {12}(753,-2)(749,-2){13}
//: {14}(755,0)(755,10)(750,10){15}
//: {16}(746,10)(742,10){17}
//: {18}(748,12)(748,22)(743,22){19}
//: {20}(739,22)(735,22)(735,22)(734,22){21}
//: {22}(741,24)(741,34)(734,34){23}
//: {24}(730,34)(726,34)(726,34)(726,34){25}
//: {26}(732,36)(1:732,46)(727,46){27}
//: {28}(723,46)(718,46){29}
//: {30}(725,48)(725,58)(718,58){31}
//: {32}(714,58)(710,58)(710,58)(710,58){33}
//: {34}(716,60)(716,70)(710,70){35}
//: {36}(706,70)(703,70)(703,70)(703,70){37}
//: {38}(708,72)(708,81)(703,81){39}
//: {40}(699,81)(694,81)(694,81)(694,81){41}
//: {42}(701,83)(701,90)(687,90){43}
//: {44}(271,818)(271,936)(-50,936)(-50,1055){45}
//: {46}(-48,1057)(-36,1057){47}
//: {48}(-52,1057)(-59,1057){49}
wire w254;    //: /sn:0 {0}(989,2260)(982,2260){1}
wire w157;    //: /sn:0 {0}(991,1821)(984,1821){1}
wire w102;    //: /sn:0 {0}(602,1672)(595,1672){1}
wire w43;    //: /sn:0 {0}(536,1671)(531,1671){1}
wire w58;    //: /sn:0 {0}(941,1944)(933,1944){1}
//: {2}(931,1942)(931,1885)(1312,1885)(1312,1066){3}
//: {4}(1312,1062)(1312,615)(582,615)(582,482)(592,482){5}
//: {6}(1310,1064)(1197,1064){7}
//: {8}(929,1944)(918,1944){9}
wire w28;    //: /sn:0 {0}(-425,1051)(-435,1051)(-435,1051)(-436,1051){1}
//: {2}(-438,1049)(-438,1005){3}
//: {4}(-438,1001)(-438,905)(259,905)(259,758){5}
//: {6}(261,756)(283,756)(283,756)(547,756){7}
//: {8}(259,754)(259,684)(125,684)(125,-219)(618,-219)(618,-70)(610,-70)(610,-60){9}
//: {10}(608,-58)(607,-58){11}
//: {12}(610,-56)(610,-48){13}
//: {14}(608,-46)(601,-46)(601,-46)(607,-46){15}
//: {16}(610,-44)(610,-35){17}
//: {18}(608,-33)(601,-33)(601,-33)(607,-33){19}
//: {20}(610,-31)(610,-22){21}
//: {22}(608,-20)(601,-20)(601,-20)(607,-20){23}
//: {24}(610,-18)(610,-9)(610,-9)(610,-9){25}
//: {26}(608,-7)(601,-7)(601,-7)(607,-7){27}
//: {28}(610,-5)(610,3){29}
//: {30}(608,5)(601,5)(601,5)(607,5){31}
//: {32}(610,7)(610,16){33}
//: {34}(608,18)(601,18)(601,18)(607,18){35}
//: {36}(610,20)(610,28){37}
//: {38}(608,30)(601,30)(601,30)(607,30){39}
//: {40}(610,32)(610,40){41}
//: {42}(608,42)(601,42)(601,42)(607,42){43}
//: {44}(610,44)(610,53){45}
//: {46}(608,55)(601,55)(601,55)(607,55){47}
//: {48}(610,57)(610,68)(607,68){49}
//: {50}(-440,1003)(-545,1003)(-545,992){51}
//: {52}(-440,1051)(-447,1051){53}
wire w169;    //: /sn:0 {0}(-228,1197)(-238,1197){1}
//: {2}(-240,1195)(-240,1141)(295,1141)(295,908){3}
//: {4}(297,906)(402,906)(402,906)(547,906){5}
//: {6}(295,904)(295,700)(974,700)(974,216)(866,216){7}
//: {8}(864,214)(864,207)(864,207)(864,211){9}
//: {10}(862,216)(854,216){11}
//: {12}(852,214)(852,207)(852,207)(852,211){13}
//: {14}(850,216)(841,216){15}
//: {16}(839,214)(839,207)(839,207)(839,211){17}
//: {18}(837,216)(828,216){19}
//: {20}(826,214)(826,207)(826,207)(826,211){21}
//: {22}(824,216)(815,216)(815,216)(815,216){23}
//: {24}(813,214)(813,207)(813,207)(813,211){25}
//: {26}(811,216)(803,216){27}
//: {28}(801,214)(801,207)(801,207)(801,211){29}
//: {30}(799,216)(790,216){31}
//: {32}(788,214)(788,207)(788,207)(788,211){33}
//: {34}(786,216)(778,216){35}
//: {36}(776,214)(776,207)(776,207)(776,211){37}
//: {38}(774,216)(766,216){39}
//: {40}(764,214)(764,207)(764,207)(764,211){41}
//: {42}(762,216)(753,216){43}
//: {44}(751,214)(751,207)(751,207)(751,211){45}
//: {46}(749,216)(738,216)(738,211){47}
//: {48}(-242,1197)(-252,1197){49}
wire w307;    //: /sn:0 {0}(13,1224)(6,1224){1}
wire w321;    //: /sn:0 {0}(-54,1662)(-61,1662){1}
wire w385;    //: /sn:0 {0}(210,1374)(203,1374){1}
wire w184;    //: /sn:0 {0}(1252,1825)(1245,1825){1}
wire w132;    //: /sn:0 {0}(553,1791)(545,1791){1}
//: {2}(543,1789)(543,1723)(1272,1723)(1272,886){3}
//: {4}(1272,882)(1272,657)(1025,657)(1025,134)(873,134)(873,131){5}
//: {6}(1270,884)(1197,884){7}
//: {8}(541,1791)(531,1791){9}
wire w269;    //: /sn:0 {0}(-315,1658)(-322,1658){1}
wire w377;    //: /sn:0 {0}(274,1085)(267,1085){1}
wire w25;    //: /sn:0 {0}(-241,798)(-254,798){1}
//: {2}(-256,796)(-256,758)(104,758)(104,620){3}
//: {4}(104,616)(104,-229)(1058,-229)(1058,706)(526,706)(526,315){5}
//: {6}(528,313)(532,313)(532,316)(534,316){7}
//: {8}(526,311)(526,304)(528,304){9}
//: {10}(532,304)(536,304)(536,304)(540,304){11}
//: {12}(530,302)(530,292)(533,292){13}
//: {14}(537,292)(546,292){15}
//: {16}(535,290)(535,280)(539,280){17}
//: {18}(543,280)(552,280){19}
//: {20}(541,278)(541,268)(545,268){21}
//: {22}(549,268)(558,268){23}
//: {24}(547,266)(547,256)(553,256){25}
//: {26}(557,256)(564,256){27}
//: {28}(555,254)(555,244)(570,244){29}
//: {30}(102,618)(89,618)(89,618)(61,618){31}
//: {32}(-258,798)(-267,798){33}
wire w65;    //: /sn:0 {0}(1244,1949)(1256,1949){1}
//: {2}(1258,1947)(1258,1904)(1322,1904)(1322,1116){3}
//: {4}(1322,1112)(1322,605)(441,605)(441,462)(463,462){5}
//: {6}(1320,1114)(1197,1114){7}
//: {8}(1258,1951)(1258,2000)(478,2000)(478,2084)(488,2084){9}
wire w210;    //: /sn:0 {0}(601,1962)(594,1962){1}
wire w121;    //: /sn:0 {0}(-604,1118)(-625,1118)(-625,1134){1}
//: {2}(-627,1136)(-878,1136)(-878,858)(-853,858){3}
//: {4}(-625,1138)(-625,1918)(37,1918)(37,1978)(211,1978)(211,1884){5}
//: {6}(213,1882)(326,1882)(326,1872)(376,1872){7}
//: {8}(209,1882)(197,1882){9}
wire w40;    //: /sn:0 {0}(726,1794)(736,1794){1}
//: {2}(740,1794)(750,1794){3}
//: {4}(738,1792)(738,1734)(1278,1734)(1278,916){5}
//: {6}(1278,912)(1278,651)(1031,651)(1031,227)(878,227)(878,211){7}
//: {8}(1276,914)(1197,914){9}
wire w92;    //: /sn:0 {0}(731,1674)(726,1674){1}
wire w283;    //: /sn:0 {0}(31,1495)(19,1495){1}
//: {2}(17,1493)(17,1445)(359,1445)(359,1188){3}
//: {4}(361,1186)(434,1186)(434,1186)(547,1186){5}
//: {6}(359,1184)(359,643)(161,643)(161,241)(336,241){7}
//: {8}(340,241)(342,241)(342,240)(348,240){9}
//: {10}(350,242)(350,243){11}
//: {12}(352,240)(357,240)(357,238)(361,238){13}
//: {14}(363,240)(363,243)(363,243)(363,241){15}
//: {16}(365,238)(370,238)(370,235)(374,235){17}
//: {18}(376,237)(376,238)(376,238)(376,238){19}
//: {20}(378,235)(382,235)(382,232)(387,232){21}
//: {22}(389,234)(389,235){23}
//: {24}(391,232)(395,232)(395,230)(399,230){25}
//: {26}(401,232)(401,232)(401,232)(401,233){27}
//: {28}(403,230)(408,230)(408,228)(412,228){29}
//: {30}(414,230)(414,231)(414,231)(414,231){31}
//: {32}(416,228)(420,228)(420,225)(425,225){33}
//: {34}(427,227)(427,228)(427,228)(427,228){35}
//: {36}(429,225)(433,225)(433,223)(437,223){37}
//: {38}(439,225)(439,226)(439,226)(439,226){39}
//: {40}(441,223)(446,223)(446,221)(450,221){41}
//: {42}(452,223)(452,224){43}
//: {44}(452,219)(452,216)(465,216)(465,221){45}
//: {46}(338,243)(338,244)(338,244)(338,245){47}
//: {48}(15,1495)(5,1495){49}
wire w30;    //: /sn:0 {0}(-853,838)(-886,838)(-886,967)(-547,967)(-547,971){1}
wire w162;    //: /sn:0 {0}(797,1818)(792,1818){1}
wire w217;    //: /sn:0 {0}(1188,1971)(1181,1971){1}
wire w149;    //: /sn:0 {0}(-635,792)(-644,792){1}
//: {2}(-646,790)(-646,740)(92,740)(92,680){3}
//: {4}(92,676)(92,-241)(675,-241)(675,93){5}
//: {6}(673,95)(665,95){7}
//: {8}(675,97)(675,107)(671,107){9}
//: {10}(667,107)(659,107){11}
//: {12}(669,109)(669,119)(666,119){13}
//: {14}(662,119)(653,119){15}
//: {16}(664,121)(664,131)(660,131){17}
//: {18}(656,131)(647,131){19}
//: {20}(658,133)(658,143)(654,143){21}
//: {22}(650,143)(641,143){23}
//: {24}(652,145)(652,155)(646,155){25}
//: {26}(642,155)(635,155){27}
//: {28}(644,157)(1:644,167)(629,167){29}
//: {30}(90,678)(79,678)(79,678)(61,678){31}
//: {32}(-648,792)(-656,792){33}
wire w146;    //: /sn:0 {0}(-260,821)(-267,821){1}
wire w222;    //: /sn:0 {0}(1251,1972)(1244,1972){1}
wire w355;    //: /sn:0 {0}(-116,1516)(-123,1516){1}
wire w248;    //: /sn:0 {0}(1056,2116)(1051,2116){1}
wire w381;    //: /sn:0 {0}(-249,1659)(-254,1659){1}
wire w286;    //: /sn:0 {0}(98,1202)(91,1202){1}
//: {2}(89,1200)(89,1163)(305,1163)(305,958){3}
//: {4}(307,956)(407,956)(407,956)(547,956){5}
//: {6}(305,954)(305,690)(984,690)(984,345)(844,345){7}
//: {8}(842,343)(842,335){9}
//: {10}(840,345)(830,345)(830,341){11}
//: {12}(830,337)(830,329){13}
//: {14}(828,339)(818,339)(818,336){15}
//: {16}(818,332)(818,323){17}
//: {18}(816,334)(806,334)(806,330){19}
//: {20}(806,326)(806,317){21}
//: {22}(804,328)(794,328)(794,324){23}
//: {24}(794,320)(794,311){25}
//: {26}(792,322)(782,322)(782,316){27}
//: {28}(782,312)(782,305){29}
//: {30}(780,314)(1:770,314)(770,308){31}
//: {32}(770,304)(770,299){33}
//: {34}(768,306)(758,306)(758,306){35}
//: {36}(758,302)(758,294){37}
//: {38}(756,304)(746,304)(746,300){39}
//: {40}(746,296)(746,288){41}
//: {42}(744,298)(734,298)(734,295){43}
//: {44}(734,291)(734,282){45}
//: {46}(732,293)(722,293)(722,276){47}
//: {48}(87,1202)(74,1202){49}
wire w173;    //: /sn:0 {0}(-101,1199)(-110,1199){1}
//: {2}(-112,1197)(-112,1150)(299,1150)(299,928){3}
//: {4}(301,926)(404,926)(404,926)(547,926){5}
//: {6}(299,924)(299,696)(978,696)(978,272)(862,272)(862,268){7}
//: {8}(862,264)(862,258)(862,258)(862,262){9}
//: {10}(860,266)(856,266)(856,263)(852,263){11}
//: {12}(850,261)(850,255)(850,255)(850,259){13}
//: {14}(848,263)(843,263)(843,261)(839,261){15}
//: {16}(837,259)(837,253)(837,253)(837,257){17}
//: {18}(835,261)(830,261)(830,259)(826,259){19}
//: {20}(824,257)(824,250)(824,250)(824,254){21}
//: {22}(822,259)(813,259)(813,256)(813,256){23}
//: {24}(811,254)(811,247)(811,247)(811,251){25}
//: {26}(809,256)(805,256)(805,254)(800,254){27}
//: {28}(798,252)(798,245)(798,245)(798,249){29}
//: {30}(796,254)(791,254)(791,252)(787,252){31}
//: {32}(785,250)(785,243)(785,243)(785,247){33}
//: {34}(783,252)(779,252)(779,250)(775,250){35}
//: {36}(773,248)(773,241)(773,241)(773,245){37}
//: {38}(771,250)(767,250)(767,247)(763,247){39}
//: {40}(761,245)(761,238)(761,238)(761,242){41}
//: {42}(759,247)(754,247)(754,244)(750,244){43}
//: {44}(748,242)(748,235)(748,235)(748,239){45}
//: {46}(746,244)(735,244)(735,237){47}
//: {48}(-114,1199)(-122,1199){49}
wire w57;    //: /sn:0 {0}(876,1943)(868,1943){1}
//: {2}(866,1941)(866,1881)(1310,1881)(1310,1056){3}
//: {4}(1310,1052)(1310,617)(606,617)(606,481)(616,481){5}
//: {6}(1308,1054)(1197,1054){7}
//: {8}(864,1943)(855,1943){9}
wire w49;    //: /sn:0 {0}(1123,1680)(1118,1680){1}
wire w318;    //: /sn:0 {0}(-53,1517)(-60,1517){1}
wire w350;    //: /sn:0 {0}(209,1666)(202,1666){1}
wire w139;    //: /sn:0 {0}(-128,823)(-133,823){1}
wire [59:0] w252;    //: /sn:0 {0}(#:553,1051)(697,1051)(697,732)(-112,732)(-112,495)(#:-94,495){1}
wire w105;    //: /sn:0 {0}(-325,820)(-332,820){1}
wire w186;    //: /sn:0 {0}(-363,1342)(-372,1342){1}
//: {2}(-374,1340)(-374,1270)(319,1270)(319,1008){3}
//: {4}(321,1006)(414,1006)(414,1006)(547,1006){5}
//: {6}(319,1004)(319,675)(704,675)(704,449){7}
//: {8}(706,447)(715,447){9}
//: {10}(702,447)(700,447)(700,437){11}
//: {12}(702,435)(707,435)(707,435)(709,435){13}
//: {14}(698,435)(695,435)(695,425){15}
//: {16}(697,423)(700,423)(700,423)(703,423){17}
//: {18}(693,423)(690,423)(690,413){19}
//: {20}(692,411)(696,411)(696,411)(697,411){21}
//: {22}(688,411)(683,411)(683,401){23}
//: {24}(685,399)(691,399){25}
//: {26}(681,399)(676,399)(676,389){27}
//: {28}(678,387)(683,387)(683,387)(685,387){29}
//: {30}(674,387)(671,387)(671,377){31}
//: {32}(673,375)(676,375)(676,375)(679,375){33}
//: {34}(669,375)(666,375)(666,365){35}
//: {36}(668,363)(672,363)(672,363)(673,363){37}
//: {38}(664,363)(659,363)(659,353){39}
//: {40}(661,351)(666,351)(666,351)(667,351){41}
//: {42}(657,351)(654,351)(654,341){43}
//: {44}(656,339)(661,339){45}
//: {46}(652,339)(648,339)(648,327)(655,327){47}
//: {48}(-376,1342)(-384,1342){49}
wire w268;    //: /sn:0 {0}(663,2255)(656,2255){1}
wire w72;    //: /sn:0 {0}(1009,2092)(997,2092){1}
//: {2}(995,2090)(995,2039)(1341,2039)(1341,1196){3}
//: {4}(1341,1192)(1341,585)(242,585)(242,245)(324,245)(324,248){5}
//: {6}(1339,1194)(1197,1194){7}
//: {8}(993,2092)(983,2092){9}
wire w94;    //: /sn:0 {0}(-520,817)(-525,817){1}
wire w33;    //: /sn:0 {0}(-102,1346)(-110,1346){1}
//: {2}(-112,1344)(-112,1286)(327,1286)(327,1048){3}
//: {4}(329,1046)(418,1046)(418,1046)(547,1046){5}
//: {6}(327,1044)(327,667)(612,667)(612,469){7}
//: {8}(614,467)(615,467){9}
//: {10}(612,465)(612,461)(611,461)(611,457){11}
//: {12}(613,455)(614,455){13}
//: {14}(611,453)(611,448)(610,448)(610,444){15}
//: {16}(612,442)(615,442)(615,442)(613,442){17}
//: {18}(610,440)(610,435)(609,435)(609,431){19}
//: {20}(611,429)(612,429)(612,429)(612,429){21}
//: {22}(609,427)(609,422)(608,422)(608,418){23}
//: {24}(610,416)(611,416){25}
//: {26}(608,414)(608,410)(607,410)(607,406){27}
//: {28}(609,404)(610,404)(610,404)(610,404){29}
//: {30}(607,402)(607,397)(606,397)(606,393){31}
//: {32}(608,391)(609,391)(609,391)(609,391){33}
//: {34}(606,389)(606,385)(605,385)(605,381){35}
//: {36}(607,379)(608,379)(608,379)(608,379){37}
//: {38}(605,377)(605,373)(604,373)(604,369){39}
//: {40}(606,367)(607,367)(607,367)(607,367){41}
//: {42}(604,365)(604,360)(603,360)(603,356){43}
//: {44}(605,354)(606,354){45}
//: {46}(603,352)(603,341)(605,341){47}
//: {48}(-114,1346)(-123,1346){49}
wire w191;    //: /sn:0 {0}(926,1820)(919,1820){1}
wire w143;    //: /sn:0 {0}(-586,816)(-593,816){1}
wire w384;    //: /sn:0 {0}(-444,1656)(-449,1656){1}
wire w107;    //: /sn:0 {0}(1057,1679)(1052,1679){1}
wire w219;    //: /sn:0 {0}(-449,1633)(-438,1633){1}
//: {2}(-434,1633)(-427,1633){3}
//: {4}(-436,1631)(-436,1561)(374,1561)(374,1238){5}
//: {6}(376,1236)(441,1236)(441,1236)(547,1236){7}
//: {8}(374,1234)(374,629)(176,629)(176,116)(337,116){9}
//: {10}(341,116)(345,116)(345,120)(349,120){11}
//: {12}(351,122)(351,127)(351,127)(351,123){13}
//: {14}(353,120)(358,120)(358,123)(362,123){15}
//: {16}(364,125)(364,130)(364,130)(364,126){17}
//: {18}(366,123)(371,123)(371,126)(375,126){19}
//: {20}(377,128)(377,135)(377,135)(377,131){21}
//: {22}(379,126)(388,126)(388,130)(388,130){23}
//: {24}(390,132)(390,139)(390,139)(390,135){25}
//: {26}(392,130)(396,130)(396,133)(401,133){27}
//: {28}(403,135)(403,142)(403,142)(403,138){29}
//: {30}(405,133)(410,133)(410,136)(414,136){31}
//: {32}(416,138)(416,145)(416,145)(416,141){33}
//: {34}(418,136)(422,136)(422,139)(426,139){35}
//: {36}(428,141)(428,148)(428,148)(428,144){37}
//: {38}(430,139)(434,139)(434,144)(438,144){39}
//: {40}(440,146)(440,153)(440,153)(440,149){41}
//: {42}(442,144)(447,144)(447,148)(451,148){43}
//: {44}(453,150)(453,157)(453,157)(453,153){45}
//: {46}(455,148)(466,148)(466,156){47}
//: {48}(339,118)(339,119){49}
wire w79;    //: /sn:0 {0}(1139,2094)(1132,2094){1}
//: {2}(1130,2092)(1130,2051)(1345,2051)(1345,1216){3}
//: {4}(1345,1212)(1345,581)(238,581)(238,184)(322,184)(322,195){5}
//: {6}(1343,1214)(1197,1214){7}
//: {8}(1128,2094)(1117,2094){9}
wire w145;    //: /sn:0 {0}(-649,815)(-656,815){1}
wire w9;    //: /sn:0 {0}(726,1651)(737,1651){1}
//: {2}(741,1651)(750,1651){3}
//: {4}(739,1649)(739,1520)(1250,1520)(1250,796){5}
//: {6}(1250,792)(1250,683)(1015,683)(1015,-183)(711,-183)(711,-70)(687,-70){7}
//: {8}(1248,794)(1197,794){9}
wire w201;    //: /sn:0 {0}(-426,1488)(-435,1488){1}
//: {2}(-437,1486)(-437,1409)(345,1409)(345,1118){3}
//: {4}(347,1116)(427,1116)(427,1116)(547,1116){5}
//: {6}(345,1114)(345,653)(319,653)(319,432)(430,432){7}
//: {8}(434,432)(437,432){9}
//: {10}(432,430)(432,420)(437,420){11}
//: {12}(441,420)(444,420){13}
//: {14}(439,418)(439,408)(444,408){15}
//: {16}(448,408)(452,408){17}
//: {18}(446,406)(446,396)(451,396){19}
//: {20}(455,396)(459,396){21}
//: {22}(453,394)(453,384)(458,384){23}
//: {24}(462,384)(466,384)(466,384)(467,384){25}
//: {26}(460,382)(460,372)(467,372){27}
//: {28}(471,372)(475,372)(475,372)(475,372){29}
//: {30}(469,370)(1:469,360)(474,360){31}
//: {32}(478,360)(483,360){33}
//: {34}(476,358)(476,348)(483,348){35}
//: {36}(487,348)(491,348)(491,348)(491,348){37}
//: {38}(485,346)(485,336)(491,336){39}
//: {40}(495,336)(498,336)(498,336)(498,336){41}
//: {42}(493,334)(493,325)(498,325){43}
//: {44}(502,325)(507,325)(507,325)(507,325){45}
//: {46}(500,323)(500,316)(514,316){47}
//: {48}(-439,1488)(-448,1488){49}
wire w55;    //: /sn:0 {0}(749,1941)(739,1941){1}
//: {2}(737,1939)(737,1873)(1306,1873)(1306,1037){3}
//: {4}(1306,1033)(1306,621)(658,621)(658,479)(668,479){5}
//: {6}(1304,1035)(1286,1035)(1286,1034)(1197,1034){7}
//: {8}(735,1941)(725,1941){9}
wire w39;    //: /sn:0 {0}(797,1675)(792,1675){1}
wire w232;    //: /sn:0 {0}(796,2112)(791,2112){1}
wire w166;    //: /sn:0 {0}(-567,793)(-580,793){1}
//: {2}(-582,791)(-582,743)(94,743)(94,670){3}
//: {4}(94,666)(94,-239)(1068,-239)(1068,169)(714,169){5}
//: {6}(712,167)(712,154){7}
//: {8}(710,169)(702,169){9}
//: {10}(700,167)(700,162)(700,162)(700,160){11}
//: {12}(700,171)(700,174)(690,174){13}
//: {14}(688,172)(688,169)(688,169)(688,166){15}
//: {16}(688,176)(688,179)(678,179){17}
//: {18}(676,177)(676,173)(676,173)(676,172){19}
//: {20}(676,181)(676,186)(666,186){21}
//: {22}(664,184)(664,179)(664,179)(664,178){23}
//: {24}(664,188)(664,191)(654,191){25}
//: {26}(652,189)(652,184){27}
//: {28}(652,193)(652,197)(640,197)(640,190){29}
//: {30}(92,668)(72,668)(72,668)(61,668){31}
//: {32}(-584,793)(-593,793){33}
wire w134;    //: /sn:0 {0}(-362,1052)(-372,1052){1}
//: {2}(-374,1050)(-374,918)(261,918)(261,768){3}
//: {4}(263,766)(286,766)(286,766)(547,766){5}
//: {6}(261,764)(261,682)(127,682)(127,-217)(645,-217)(645,-70)(638,-70)(638,-60){7}
//: {8}(636,-58)(629,-58)(629,-58)(633,-58){9}
//: {10}(638,-56)(638,-52)(636,-52)(636,-48){11}
//: {12}(634,-46)(627,-46)(627,-46)(631,-46){13}
//: {14}(636,-44)(636,-39)(635,-39)(635,-35){15}
//: {16}(633,-33)(630,-33){17}
//: {18}(635,-31)(635,-26)(633,-26)(633,-22){19}
//: {20}(631,-20)(624,-20)(624,-20)(628,-20){21}
//: {22}(633,-18)(633,-9)(632,-9)(632,-9){23}
//: {24}(630,-7)(623,-7)(623,-7)(627,-7){25}
//: {26}(632,-5)(632,-1)(631,-1)(631,4){27}
//: {28}(629,6)(622,6)(622,6)(626,6){29}
//: {30}(631,8)(631,13)(630,13)(630,17){31}
//: {32}(628,19)(621,19)(621,19)(625,19){33}
//: {34}(630,21)(630,25)(629,25)(629,29){35}
//: {36}(627,31)(620,31)(620,31)(624,31){37}
//: {38}(629,33)(629,37)(628,37)(628,41){39}
//: {40}(626,43)(619,43)(619,43)(623,43){41}
//: {42}(628,45)(628,50)(626,50)(626,54){43}
//: {44}(624,56)(617,56)(617,56)(621,56){45}
//: {46}(626,58)(626,69)(620,69){47}
//: {48}(-376,1052)(-383,1052){49}
wire w214;    //: /sn:0 {0}(730,1964)(725,1964){1}
wire w141;    //: /sn:0 {0}(547,1326)(450,1326)(450,1326)(394,1326){1}
//: {2}(392,1324)(392,611)(194,611)(194,-155)(537,-155)(537,-57){3}
//: {4}(535,-55)(534,-55)(534,-55)(533,-55){5}
//: {6}(537,-53)(537,-51)(539,-51)(539,-45){7}
//: {8}(541,-43)(551,-43)(551,-43)(537,-43){9}
//: {10}(539,-41)(539,-36)(543,-36)(543,-32){11}
//: {12}(541,-30)(538,-30)(538,-30)(540,-30){13}
//: {14}(543,-28)(543,-23)(547,-23)(547,-19){15}
//: {16}(545,-17)(544,-17)(544,-17)(544,-17){17}
//: {18}(547,-15)(547,-11)(551,-11)(551,-6){19}
//: {20}(549,-4)(548,-4){21}
//: {22}(551,-2)(551,2)(554,2)(554,6){23}
//: {24}(552,8)(552,8)(552,8)(551,8){25}
//: {26}(554,10)(554,15)(558,15)(558,18){27}
//: {28}(556,20)(555,20)(555,20)(555,20){29}
//: {30}(558,22)(558,26)(562,26)(562,31){31}
//: {32}(560,33)(559,33)(559,33)(559,33){33}
//: {34}(562,35)(562,39)(565,39)(565,43){35}
//: {36}(563,45)(562,45)(562,45)(562,45){37}
//: {38}(565,47)(565,52)(569,52)(569,56){39}
//: {40}(567,58)(566,58){41}
//: {42}(571,58)(574,58)(574,71)(570,71){43}
//: {44}(392,1328)(392,1609)(148,1609)(148,1640){45}
//: {46}(150,1642)(160,1642){47}
//: {48}(146,1642)(138,1642){49}
wire w386;    //: /sn:0 {0}(210,1521)(203,1521){1}
wire w14;    //: /sn:0 {0}(1197,824)(1254,824){1}
//: {2}(1256,822)(1256,677)(1009,677)(1009,-39)(773,-39){3}
//: {4}(1256,826)(1256,1531)(928,1531)(928,1652){5}
//: {6}(930,1654)(942,1654){7}
//: {8}(926,1654)(919,1654){9}
wire w220;    //: /sn:0 {0}(1122,1970)(1117,1970){1}
wire [5:0] w38;    //: /sn:0 {0}(297,12)(297,18)(#:29,18)(29,493)(#:3,493){1}
wire w250;    //: /sn:0 {0}(535,2108)(530,2108){1}
wire w292;    //: /sn:0 {0}(145,1226)(140,1226){1}
wire w181;    //: /sn:0 {0}(225,1204)(218,1204){1}
//: {2}(216,1202)(216,1171)(309,1171)(309,978){3}
//: {4}(311,976)(409,976)(409,976)(547,976){5}
//: {6}(309,974)(309,686)(988,686)(988,401)(816,401){7}
//: {8}(814,399)(814,397){9}
//: {10}(812,401)(803,401)(803,394){11}
//: {12}(803,390)(803,388)(803,388)(803,388){13}
//: {14}(801,392)(792,392)(792,386){15}
//: {16}(792,382)(792,379)(792,379)(792,379){17}
//: {18}(790,384)(781,384)(781,378){19}
//: {20}(781,374)(781,370)(781,370)(781,370){21}
//: {22}(779,376)(770,376)(770,368){23}
//: {24}(770,364)(770,361)(770,361)(770,361){25}
//: {26}(768,366)(759,366)(759,358){27}
//: {28}(759,354)(759,352)(759,352)(759,352){29}
//: {30}(1:757,356)(748,356)(748,349){31}
//: {32}(748,345)(748,343)(748,343)(748,343){33}
//: {34}(746,347)(737,347)(737,340){35}
//: {36}(737,336)(737,334)(737,334)(737,334){37}
//: {38}(735,338)(726,338)(726,334){39}
//: {40}(726,330)(726,326)(726,326)(726,325){41}
//: {42}(724,332)(715,332)(715,323){43}
//: {44}(715,319)(715,316)(715,316)(715,316){45}
//: {46}(713,321)(705,321)(705,307){47}
//: {48}(214,1204)(204,1204){49}
wire w302;    //: /sn:0 {0}(-116,1369)(-123,1369){1}
wire w3;    //: /sn:0 {0}(616,1649)(606,1649){1}
//: {2}(604,1647)(604,1512)(1246,1512)(1246,776){3}
//: {4}(1246,772)(1246,687)(1019,687)(1019,-187)(640,-187)(640,-72)(635,-72){5}
//: {6}(1244,774)(1197,774){7}
//: {8}(602,1649)(595,1649){9}
wire w204;    //: /sn:0 {0}(-229,1491)(-241,1491){1}
//: {2}(-243,1489)(-243,1425)(351,1425)(351,1148){3}
//: {4}(353,1146)(430,1146)(430,1146)(547,1146){5}
//: {6}(351,1144)(351,489)(285,489)(285,346)(366,346){7}
//: {8}(368,344)(368,338)(377,338){9}
//: {10}(379,340)(379,342)(379,342)(379,344){11}
//: {12}(379,336)(379,330)(388,330){13}
//: {14}(390,332)(390,334)(390,334)(390,336){15}
//: {16}(390,328)(390,321)(400,321){17}
//: {18}(402,323)(402,330)(402,330)(402,329){19}
//: {20}(402,319)(402,312)(412,312){21}
//: {22}(414,314)(414,320)(414,320)(414,321){23}
//: {24}(414,310)(414,306)(423,306){25}
//: {26}(425,308)(425,313)(425,313)(425,313){27}
//: {28}(425,304)(425,299)(435,299){29}
//: {30}(437,301)(437,305)(437,305)(437,305){31}
//: {32}(437,297)(437,293)(447,293){33}
//: {34}(449,295)(449,298)(449,298)(449,297){35}
//: {36}(449,291)(449,286)(459,286){37}
//: {38}(461,288)(461,290)(461,290)(461,290){39}
//: {40}(461,284)(461,277)(471,277){41}
//: {42}(473,279)(473,281)(473,281)(473,282){43}
//: {44}(473,275)(473,272)(485,272)(485,275){45}
//: {46}(368,348)(368,351)(368,351)(368,352){47}
//: {48}(-245,1491)(-253,1491){49}
wire w75;    //: /sn:0 {0}(791,2089)(808,2089){1}
//: {2}(812,2089)(813,2089){3}
//: {4}(810,2087)(810,2023)(1335,2023)(1335,1166){5}
//: {6}(1335,1162)(1335,591)(248,591)(248,317)(344,317)(344,327){7}
//: {8}(1333,1164)(1197,1164){9}
wire w360;    //: /sn:0 {0}(96,1641)(87,1641){1}
//: {2}(85,1639)(85,1605)(390,1605)(390,1318){3}
//: {4}(392,1316)(449,1316)(449,1316)(547,1316){5}
//: {6}(390,1314)(390,613)(192,613)(192,-153)(511,-153)(511,-51){7}
//: {8}(509,-49)(508,-49)(508,-49)(507,-49){9}
//: {10}(511,-47)(511,-45)(515,-45)(515,-40){11}
//: {12}(513,-38)(512,-38){13}
//: {14}(515,-36)(515,-31)(520,-31)(520,-27){15}
//: {16}(518,-25)(515,-25)(515,-25)(517,-25){17}
//: {18}(520,-23)(520,-18)(526,-18)(526,-14){19}
//: {20}(524,-12)(523,-12)(523,-12)(523,-12){21}
//: {22}(526,-10)(526,-6)(531,-6)(531,-2){23}
//: {24}(529,0)(528,0){25}
//: {26}(531,2)(531,6)(536,6)(536,10){27}
//: {28}(534,12)(534,12)(534,12)(533,12){29}
//: {30}(536,14)(536,19)(541,19)(541,23){31}
//: {32}(539,25)(538,25)(538,25)(538,25){33}
//: {34}(541,27)(541,31)(546,31)(546,35){35}
//: {36}(544,37)(543,37)(543,37)(543,37){37}
//: {38}(546,39)(546,43)(551,43)(551,47){39}
//: {40}(549,49)(548,49)(548,49)(548,49){41}
//: {42}(551,51)(551,56)(556,56)(556,60){43}
//: {44}(554,62)(553,62){45}
//: {46}(558,62)(561,62)(561,75)(558,75){47}
//: {48}(83,1641)(72,1641){49}
wire w379;    //: /sn:0 {0}(-181,1078)(-186,1078){1}
wire w276;    //: /sn:0 {0}(924,2259)(917,2259){1}
wire w215;    //: /sn:0 {0}(224,1498)(215,1498){1}
//: {2}(213,1496)(213,1462)(365,1462)(365,1218){3}
//: {4}(367,1216)(437,1216)(437,1216)(547,1216){5}
//: {6}(365,1214)(365,637)(167,637)(167,164)(335,164){7}
//: {8}(339,164)(343,164)(343,166)(347,166){9}
//: {10}(349,168)(349,175)(349,175)(349,171){11}
//: {12}(351,166)(356,166)(356,167)(360,167){13}
//: {14}(362,169)(362,176)(362,176)(362,172){15}
//: {16}(364,167)(369,167)(369,169)(373,169){17}
//: {18}(375,171)(375,178)(375,178)(375,174){19}
//: {20}(377,169)(386,169)(386,170)(386,170){21}
//: {22}(388,172)(388,179)(388,179)(388,175){23}
//: {24}(390,170)(394,170)(394,171)(399,171){25}
//: {26}(401,173)(401,180)(401,180)(401,176){27}
//: {28}(403,171)(408,171)(408,172)(412,172){29}
//: {30}(414,174)(414,181)(414,181)(414,177){31}
//: {32}(416,172)(420,172)(420,173)(424,173){33}
//: {34}(426,175)(426,182)(426,182)(426,178){35}
//: {36}(428,173)(432,173)(432,174)(436,174){37}
//: {38}(438,176)(438,183)(438,183)(438,179){39}
//: {40}(440,174)(445,174)(445,176)(449,176){41}
//: {42}(451,178)(451,185)(451,185)(451,181){43}
//: {44}(453,176)(464,176)(464,182){45}
//: {46}(337,166)(337,173)(337,173)(337,169){47}
//: {48}(211,1498)(203,1498){49}
wire w311;    //: /sn:0 {0}(-182,1515)(-187,1515){1}
wire w156;    //: /sn:0 {0}(1197,904)(1274,904){1}
//: {2}(1276,902)(1276,653)(1029,653)(1029,192)(878,192)(878,187){3}
//: {4}(1276,906)(1276,1730)(671,1730)(671,1791){5}
//: {6}(673,1793)(684,1793){7}
//: {8}(669,1793)(658,1793){9}
wire w41;    //: /sn:0 {0}(-309,797)(-319,797){1}
//: {2}(-321,795)(-321,755)(102,755)(102,630){3}
//: {4}(102,626)(102,-231)(1060,-231)(1060,708)(586,708)(586,331){5}
//: {6}(588,329)(592,329){7}
//: {8}(586,327)(586,319){9}
//: {10}(588,317)(595,317)(595,317)(592,317){11}
//: {12}(586,315)(586,306){13}
//: {14}(588,304)(592,304){15}
//: {16}(586,302)(586,294){17}
//: {18}(588,292)(590,292)(590,292)(592,292){19}
//: {20}(586,290)(586,282){21}
//: {22}(588,280)(590,280)(590,280)(592,280){23}
//: {24}(586,278)(586,269){25}
//: {26}(588,267)(592,267){27}
//: {28}(586,265)(586,254)(592,254){29}
//: {30}(100,628)(76,628)(76,628)(61,628){31}
//: {32}(-323,797)(-332,797){33}
wire [3:0] w36;    //: /sn:0 {0}(#:8,584)(25,584)(25,15)(251,15)(251,12){1}
wire w324;    //: /sn:0 {0}(211,1084)(204,1084){1}
wire w242;    //: /sn:0 {0}(1188,2118)(1181,2118){1}
wire w82;    //: /sn:0 {0}(529,2230)(540,2230){1}
//: {2}(544,2230)(551,2230){3}
//: {4}(542,2228)(542,2159)(1354,2159)(1354,1246){5}
//: {6}(1354,1242)(1354,570)(205,570)(205,112)(325,112)(325,115){7}
//: {8}(1352,1244)(1197,1244){9}
wire w74;    //: /sn:0 {0}(876,2090)(863,2090){1}
//: {2}(861,2088)(861,2028)(1337,2028)(1337,1176){3}
//: {4}(1337,1172)(1337,589)(246,589)(246,296)(333,296)(333,301){5}
//: {6}(1335,1174)(1197,1174){7}
//: {8}(859,2090)(855,2090){9}
wire w35;    //: /sn:0 {0}(-165,1345)(-176,1345){1}
//: {2}(-178,1343)(-178,1282)(325,1282)(325,1038){3}
//: {4}(327,1036)(417,1036)(417,1036)(547,1036){5}
//: {6}(325,1034)(325,669)(637,669)(637,469){7}
//: {8}(639,467)(640,467)(640,467)(641,467){9}
//: {10}(637,465)(637,463)(636,463)(636,457){11}
//: {12}(638,455)(639,455){13}
//: {14}(636,453)(636,448)(634,448)(634,444){15}
//: {16}(636,442)(639,442)(639,442)(637,442){17}
//: {18}(634,440)(634,435)(631,435)(631,431){19}
//: {20}(633,429)(634,429)(634,429)(634,429){21}
//: {22}(631,427)(631,423)(628,423)(628,418){23}
//: {24}(630,416)(631,416){25}
//: {26}(628,414)(628,410)(626,410)(626,406){27}
//: {28}(628,404)(629,404){29}
//: {30}(626,402)(626,397)(624,397)(624,393){31}
//: {32}(626,391)(627,391)(627,391)(627,391){33}
//: {34}(624,389)(624,385)(621,385)(621,380){35}
//: {36}(623,378)(624,378)(624,378)(624,378){37}
//: {38}(621,376)(621,372)(619,372)(619,368){39}
//: {40}(621,366)(622,366)(622,366)(622,366){41}
//: {42}(619,364)(619,359)(617,359)(617,355){43}
//: {44}(619,353)(620,353){45}
//: {46}(615,353)(612,353)(612,340)(617,340){47}
//: {48}(-180,1345)(-187,1345){49}
wire w91;    //: /sn:0 {0}(854,2235)(863,2235){1}
//: {2}(867,2235)(875,2235){3}
//: {4}(865,2233)(865,2186)(1364,2186)(1364,1296){5}
//: {6}(1364,1292)(1364,560)(215,560)(215,-166)(412,-166)(412,-22)(406,-22){7}
//: {8}(1362,1294)(1197,1294){9}
wire [5:0] w101;    //: /sn:0 {0}(#:343,12)(343,20)(33,20)(33,538)(3,538){1}
wire w163;    //: /sn:0 {0}(-294,1053)(-309,1053){1}
//: {2}(-311,1051)(-311,921)(263,921)(263,778){3}
//: {4}(265,776)(290,776)(290,776)(547,776){5}
//: {6}(263,774)(263,680)(129,680)(129,-215)(662,-215)(662,-60){7}
//: {8}(660,-58)(654,-58)(654,-58)(658,-58){9}
//: {10}(662,-56)(662,-52)(659,-52)(659,-48){11}
//: {12}(657,-46)(655,-46){13}
//: {14}(659,-44)(659,-39)(657,-39)(657,-35){15}
//: {16}(655,-33)(649,-33)(649,-33)(653,-33){17}
//: {18}(657,-31)(657,-26)(655,-26)(655,-22){19}
//: {20}(653,-20)(646,-20)(646,-20)(650,-20){21}
//: {22}(655,-18)(655,-9)(652,-9)(652,-9){23}
//: {24}(650,-7)(643,-7)(643,-7)(647,-7){25}
//: {26}(652,-5)(652,-1)(650,-1)(650,4){27}
//: {28}(648,6)(641,6)(641,6)(645,6){29}
//: {30}(650,8)(650,13)(648,13)(648,17){31}
//: {32}(646,19)(639,19)(639,19)(643,19){33}
//: {34}(648,21)(648,25)(646,25)(646,29){35}
//: {36}(644,31)(637,31)(637,31)(641,31){37}
//: {38}(646,33)(646,37)(643,37)(643,41){39}
//: {40}(641,43)(634,43)(634,43)(638,43){41}
//: {42}(643,45)(643,50)(640,50)(640,54){43}
//: {44}(638,56)(631,56)(631,56)(635,56){45}
//: {46}(640,58)(640,69)(633,69){47}
//: {48}(-313,1053)(-320,1053){49}
wire w382;    //: /sn:0 {0}(12,1371)(5,1371){1}
wire w22;    //: /sn:0 {0}(649,315)(636,315){1}
//: {2}(634,313)(634,305){3}
//: {4}(636,303)(641,303)(641,303)(643,303){5}
//: {6}(632,303)(629,303)(629,293){7}
//: {8}(631,291)(634,291)(634,291)(637,291){9}
//: {10}(627,291)(624,291)(624,281){11}
//: {12}(626,279)(631,279){13}
//: {14}(622,279)(617,279)(617,269){15}
//: {16}(619,267)(625,267){17}
//: {18}(615,267)(612,267)(612,257){19}
//: {20}(614,255)(619,255){21}
//: {22}(610,255)(606,255)(606,243)(613,243){23}
//: {24}(634,317)(634,710)(1062,710)(1062,-233)(100,-233)(100,636){25}
//: {26}(98,638)(88,638)(88,638)(61,638){27}
//: {28}(100,640)(100,752)(-385,752)(-385,794){29}
//: {30}(-383,796)(-374,796){31}
//: {32}(-387,796)(-395,796){33}
wire w265;    //: /sn:0 {0}(-230,1636)(-240,1636){1}
//: {2}(-242,1634)(-242,1578)(380,1578)(380,1268){3}
//: {4}(382,1266)(444,1266)(444,1266)(547,1266){5}
//: {6}(380,1264)(380,623)(182,623)(182,24)(371,24)(371,32){7}
//: {8}(373,34)(383,34)(383,39){9}
//: {10}(383,43)(383,46){11}
//: {12}(385,41)(395,41)(395,46){13}
//: {14}(395,50)(395,54){15}
//: {16}(397,48)(407,48)(407,53){17}
//: {18}(407,57)(407,61){19}
//: {20}(409,55)(419,55)(419,60){21}
//: {22}(419,64)(419,68)(419,68)(419,69){23}
//: {24}(421,62)(431,62)(431,69){25}
//: {26}(431,73)(431,77)(431,77)(431,77){27}
//: {28}(433,71)(1:443,71)(443,76){29}
//: {30}(443,80)(443,85){31}
//: {32}(445,78)(455,78)(455,85){33}
//: {34}(455,89)(455,93)(455,93)(455,93){35}
//: {36}(457,87)(467,87)(467,93){37}
//: {38}(467,97)(467,100)(467,100)(467,100){39}
//: {40}(469,95)(478,95)(478,100){41}
//: {42}(480,102)(487,102)(487,116){43}
//: {44}(478,104)(478,109)(478,109)(478,109){45}
//: {46}(371,36)(371,39){47}
//: {48}(-244,1636)(-254,1636){49}
wire w296;    //: /sn:0 {0}(-61,1639)(-53,1639){1}
//: {2}(-49,1639)(-38,1639){3}
//: {4}(-51,1637)(-51,1595)(386,1595)(386,1298){5}
//: {6}(388,1296)(447,1296)(447,1296)(547,1296){7}
//: {8}(386,1294)(386,617)(188,617)(188,-149)(457,-149)(457,-32){9}
//: {10}(459,-30)(465,-30)(465,-21){11}
//: {12}(463,-19)(461,-19)(461,-19)(459,-19){13}
//: {14}(467,-19)(473,-19)(473,-10){15}
//: {16}(471,-8)(469,-8)(469,-8)(467,-8){17}
//: {18}(475,-8)(482,-8)(482,2){19}
//: {20}(480,4)(473,4)(473,4)(474,4){21}
//: {22}(484,4)(491,4)(491,14){23}
//: {24}(489,16)(483,16)(483,16)(482,16){25}
//: {26}(493,16)(497,16)(497,25){27}
//: {28}(495,27)(490,27)(490,27)(490,27){29}
//: {30}(499,27)(504,27)(504,37){31}
//: {32}(502,39)(498,39)(498,39)(498,39){33}
//: {34}(506,39)(510,39)(510,49){35}
//: {36}(508,51)(505,51)(505,51)(506,51){37}
//: {38}(512,51)(517,51)(517,61){39}
//: {40}(515,63)(513,63)(513,63)(513,63){41}
//: {42}(519,63)(526,63)(526,73){43}
//: {44}(524,75)(522,75)(522,75)(521,75){45}
//: {46}(528,75)(531,75)(531,87)(528,87){47}
//: {48}(455,-30)(452,-30)(452,-30)(451,-30){49}
wire w332;    //: /sn:0 {0}(162,1060)(150,1060){1}
//: {2}(148,1058)(148,949)(277,949)(277,848){3}
//: {4}(279,846)(328,846)(328,846)(547,846){5}
//: {6}(277,844)(277,666)(143,666)(143,-201)(998,-201)(998,60)(835,60){7}
//: {8}(833,58)(833,55)(833,55)(833,54){9}
//: {10}(833,62)(833,68)(824,68){11}
//: {12}(822,66)(822,64)(822,64)(822,62){13}
//: {14}(822,70)(822,76)(813,76){15}
//: {16}(811,74)(811,72)(811,72)(811,70){17}
//: {18}(811,78)(811,85)(801,85){19}
//: {20}(799,83)(799,76)(799,76)(799,77){21}
//: {22}(799,87)(799,94)(789,94){23}
//: {24}(787,92)(787,86)(787,86)(787,85){25}
//: {26}(787,96)(787,100)(778,100){27}
//: {28}(776,98)(776,93)(776,93)(776,93){29}
//: {30}(776,102)(776,107)(766,107){31}
//: {32}(764,105)(764,101)(764,101)(764,101){33}
//: {34}(764,109)(764,113)(754,113){35}
//: {36}(752,111)(752,108)(752,108)(752,109){37}
//: {38}(752,115)(752,120)(742,120){39}
//: {40}(740,118)(740,116)(740,116)(740,116){41}
//: {42}(740,122)(740,129)(730,129){43}
//: {44}(728,127)(728,125)(728,125)(728,124){45}
//: {46}(728,131)(728,134)(716,134)(716,131){47}
//: {48}(146,1060)(140,1060){49}
wire w172;    //: /sn:0 {0}(731,1817)(726,1817){1}
wire w228;    //: /sn:0 {0}(-188,1637)(-178,1637){1}
//: {2}(-174,1637)(-166,1637){3}
//: {4}(-176,1635)(-176,1583)(382,1583)(382,1278){5}
//: {6}(384,1276)(445,1276)(445,1276)(547,1276){7}
//: {8}(382,1274)(382,621)(184,621)(184,-145)(386,-145)(386,5){9}
//: {10}(388,7)(397,7)(397,14){11}
//: {12}(397,18)(397,20)(397,20)(397,20){13}
//: {14}(399,16)(408,16)(408,22){15}
//: {16}(408,26)(408,29)(408,29)(408,29){17}
//: {18}(410,24)(419,24)(419,30){19}
//: {20}(419,34)(419,38)(419,38)(419,38){21}
//: {22}(421,32)(430,32)(430,40){23}
//: {24}(430,44)(430,47)(430,47)(430,47){25}
//: {26}(432,42)(441,42)(441,50){27}
//: {28}(441,54)(441,56)(441,56)(441,56){29}
//: {30}(1:443,52)(452,52)(452,59){31}
//: {32}(452,63)(452,65)(452,65)(452,65){33}
//: {34}(454,61)(463,61)(463,68){35}
//: {36}(463,72)(463,74)(463,74)(463,74){37}
//: {38}(465,70)(474,70)(474,74){39}
//: {40}(474,78)(474,82)(474,82)(474,83){41}
//: {42}(476,76)(485,76)(485,85){43}
//: {44}(485,89)(485,92)(485,92)(485,92){45}
//: {46}(487,87)(495,87)(495,101){47}
//: {48}(386,9)(386,11){49}
wire w12;    //: /sn:0 {0}(1076,1656)(1064,1656){1}
//: {2}(1062,1654)(1062,1538)(1260,1538)(1260,846){3}
//: {4}(1260,842)(1260,673)(1005,673)(1005,18)(826,18)(826,11){5}
//: {6}(1258,844)(1197,844){7}
//: {8}(1060,1656)(1052,1656){9}
wire w226;    //: /sn:0 {0}(925,1967)(918,1967){1}
wire w309;    //: /sn:0 {0}(-314,1366)(-321,1366){1}
wire w78;    //: /sn:0 {0}(-454,818)(-459,818){1}
wire w200;    //: /sn:0 {0}(990,1968)(983,1968){1}
wire w365;    //: /sn:0 {0}(-183,1660)(-188,1660){1}
wire w27;    //: /sn:0 {0}(-175,799)(-185,799){1}
//: {2}(-187,797)(-187,761)(106,761)(106,610){3}
//: {4}(106,606)(106,238)(487,238){5}
//: {6}(491,238)(499,238){7}
//: {8}(501,236)(501,233)(511,233){9}
//: {10}(513,235)(513,238)(513,238)(513,241){11}
//: {12}(513,231)(513,228)(523,228){13}
//: {14}(525,230)(525,234)(525,234)(525,235){15}
//: {16}(525,226)(525,221)(535,221){17}
//: {18}(537,219)(537,216)(547,216){19}
//: {20}(549,214)(549,210)(561,210)(561,217){21}
//: {22}(549,218)(549,223){23}
//: {24}(537,223)(537,228)(537,228)(537,229){25}
//: {26}(501,240)(501,247){27}
//: {28}(489,240)(489,246)(489,246)(489,253){29}
//: {30}(104,608)(86,608)(86,608)(61,608){31}
//: {32}(-189,799)(-199,799){33}
wire w257;    //: /sn:0 {0}(795,2257)(790,2257){1}
wire w86;    //: /sn:0 {0}(614,2231)(604,2231){1}
//: {2}(602,2229)(602,2164)(1356,2164)(1356,1256){3}
//: {4}(1356,1252)(1356,568)(207,568)(207,86)(334,86)(334,89){5}
//: {6}(1354,1254)(1197,1254){7}
//: {8}(600,2231)(593,2231){9}
wire w80;    //: /sn:0 {0}(1075,2093)(1064,2093){1}
//: {2}(1062,2091)(1062,2045)(1343,2045)(1343,1206){3}
//: {4}(1343,1202)(1343,583)(240,583)(240,212)(323,212)(323,221){5}
//: {6}(1341,1204)(1197,1204){7}
//: {8}(1060,2093)(1051,2093){9}
wire w29;    //: /sn:0 {0}(-111,800)(-120,800){1}
//: {2}(-122,798)(-122,764)(108,764)(108,600){3}
//: {4}(108,596)(108,189)(473,189){5}
//: {6}(477,189)(481,189)(481,189)(485,189){7}
//: {8}(489,189)(498,189){9}
//: {10}(502,189)(510,189){11}
//: {12}(514,189)(519,189)(519,189)(523,189){13}
//: {14}(527,189)(530,189)(530,189)(535,189){15}
//: {16}(539,189)(550,189)(550,195){17}
//: {18}(537,191)(537,193)(537,193)(537,195){19}
//: {20}(525,191)(525,193)(525,193)(525,195){21}
//: {22}(512,191)(512,195){23}
//: {24}(500,191)(500,198)(500,198)(500,195){25}
//: {26}(487,191)(487,195){27}
//: {28}(475,191)(475,193)(475,193)(475,195){29}
//: {30}(106,598)(79,598)(79,598)(61,598){31}
//: {32}(-124,800)(-133,800){33}
wire w378;    //: /sn:0 {0}(-443,1364)(-448,1364){1}
wire w42;    //: /sn:0 {0}(1197,894)(1272,894){1}
//: {2}(1274,892)(1274,655)(1027,655)(1027,160)(876,160)(876,157){3}
//: {4}(1274,896)(1274,1727)(608,1727)(608,1790){5}
//: {6}(610,1792)(616,1792){7}
//: {8}(606,1792)(595,1792){9}
wire w264;    //: /sn:0 {0}(729,2256)(724,2256){1}
wire w281;    //: /sn:0 {0}(-313,1219)(-320,1219){1}
wire w370;    //: /sn:0 {0}(12,1518)(5,1518){1}
wire w317;    //: /sn:0 {0}(266,1352)(278,1352){1}
//: {2}(280,1350)(280,1312)(339,1312)(339,1108){3}
//: {4}(341,1106)(424,1106)(424,1106)(547,1106){5}
//: {6}(339,1104)(339,455)(459,455)(459,450){7}
//: {8}(461,448)(469,448){9}
//: {10}(459,446)(459,436)(463,436){11}
//: {12}(467,436)(475,436){13}
//: {14}(465,434)(465,424)(468,424){15}
//: {16}(472,424)(481,424){17}
//: {18}(470,422)(470,412)(474,412){19}
//: {20}(478,412)(487,412){21}
//: {22}(476,410)(476,400)(480,400){23}
//: {24}(484,400)(493,400){25}
//: {26}(482,398)(482,388)(488,388){27}
//: {28}(492,388)(499,388){29}
//: {30}(490,386)(1:490,376)(496,376){31}
//: {32}(500,376)(505,376){33}
//: {34}(498,374)(498,371)(500,371)(500,366){35}
//: {36}(502,364)(506,364)(506,364)(510,364){37}
//: {38}(500,362)(500,352)(504,352){39}
//: {40}(508,352)(516,352){41}
//: {42}(506,350)(506,340)(509,340){43}
//: {44}(513,340)(522,340){45}
//: {46}(511,338)(511,328)(528,328){47}
//: {48}(280,1354)(280,1403)(-500,1403)(-500,1487)(-490,1487){49}
wire w277;    //: /sn:0 {0}(78,1519)(73,1519){1}
wire w247;    //: /sn:0 {0}(1251,2119)(1244,2119){1}
wire w112;    //: /sn:0 {0}(-575,1108)(-572,1108)(-572,927)(-548,927){1}
wire w60;    //: /sn:0 {0}(1075,1946)(1067,1946){1}
//: {2}(1065,1944)(1065,1893)(1316,1893)(1316,1086){3}
//: {4}(1316,1082)(1316,611)(520,611)(520,483)(537,483){5}
//: {6}(1314,1084)(1197,1084){7}
//: {8}(1063,1946)(1051,1946){9}
wire w46;    //: /sn:0 {0}(856,1796)(864,1796){1}
//: {2}(868,1796)(877,1796){3}
//: {4}(866,1794)(866,1741)(1282,1741)(1282,936){5}
//: {6}(1282,932)(1282,647)(1035,647)(1035,268)(876,268)(876,264){7}
//: {8}(1280,934)(1197,934){9}
wire w175;    //: /sn:0 {0}(1189,1824)(1182,1824){1}
wire w336;    //: /sn:0 {0}(274,1667)(265,1667){1}
wire w15;    //: /sn:0 {0}(877,1653)(867,1653){1}
//: {2}(865,1651)(865,1528)(1254,1528)(1254,816){3}
//: {4}(1254,812)(1254,679)(1011,679)(1011,-51)(737,-51){5}
//: {6}(1252,814)(1197,814){7}
//: {8}(863,1653)(856,1653){9}
wire w291;    //: /sn:0 {0}(-117,1661)(-124,1661){1}
wire w109;    //: /sn:0 {0}(-762,790)(-808,790)(-808,791)(-855,791){1}
wire w129;    //: /sn:0 {0}(-194,822)(-199,822){1}
wire w306;    //: /sn:0 {0}(273,1375)(266,1375){1}
wire w114;    //: /sn:0 {0}(271,1802)(271,1719)(271,1719)(271,1796){1}
wire w97;    //: /sn:0 {0}(1074,2238)(1065,2238){1}
//: {2}(1063,2236)(1063,2201)(1370,2201)(1370,1326){3}
//: {4}(1370,1322)(1370,554)(221,554)(221,-172)(508,-172)(508,-63)(502,-63){5}
//: {6}(1368,1324)(1197,1324){7}
//: {8}(1061,2238)(1050,2238){9}
wire w229;    //: /sn:0 {0}(990,2115)(983,2115){1}
wire w331;    //: /sn:0 {0}(-181,1221)(-186,1221){1}
wire w64;    //: /sn:0 {0}(265,1644)(276,1644){1}
//: {2}(278,1642)(278,1620)(396,1620)(396,1348){3}
//: {4}(398,1346)(452,1346)(452,1346)(547,1346){5}
//: {6}(396,1344)(396,607)(198,607)(198,-159)(587,-159)(587,-60){7}
//: {8}(585,-58)(584,-58){9}
//: {10}(587,-56)(587,-52)(588,-52)(588,-48){11}
//: {12}(586,-46)(585,-46){13}
//: {14}(588,-44)(588,-39)(589,-39)(589,-35){15}
//: {16}(587,-33)(584,-33)(584,-33)(586,-33){17}
//: {18}(589,-31)(589,-26)(590,-26)(590,-22){19}
//: {20}(588,-20)(587,-20)(587,-20)(587,-20){21}
//: {22}(590,-18)(590,-13)(591,-13)(591,-9){23}
//: {24}(589,-7)(588,-7){25}
//: {26}(591,-5)(591,-1)(592,-1)(592,3){27}
//: {28}(590,5)(589,5)(589,5)(589,5){29}
//: {30}(592,7)(592,12)(593,12)(593,16){31}
//: {32}(591,18)(590,18)(590,18)(590,18){33}
//: {34}(593,20)(593,24)(594,24)(594,28){35}
//: {36}(592,30)(591,30)(591,30)(591,30){37}
//: {38}(594,32)(594,36)(595,36)(595,40){39}
//: {40}(593,42)(592,42)(592,42)(592,42){41}
//: {42}(595,44)(595,49)(596,49)(596,53){43}
//: {44}(594,55)(593,55){45}
//: {46}(596,57)(596,68)(594,68){47}
//: {48}(278,1646)(278,1656)(294,1656)(294,1697)(-651,1697)(-651,1191){49}
wire w245;    //: /sn:0 {0}(1122,2117)(1117,2117){1}
wire w267;    //: /sn:0 {0}(1187,2263)(1180,2263){1}
wire w261;    //: /sn:0 {0}(-378,1657)(-385,1657){1}
wire w285;    //: /sn:0 {0}(-248,1514)(-253,1514){1}
wire w63;    //: /sn:0 {0}(1202,1948)(1199,1948){1}
//: {2}(1197,1946)(1197,1901)(1320,1901)(1320,1106){3}
//: {4}(1320,1102)(1320,607)(469,607)(469,471)(488,471){5}
//: {6}(1318,1104)(1197,1104){7}
//: {8}(1195,1948)(1181,1948){9}
wire w361;    //: /sn:0 {0}(77,1664)(72,1664){1}
wire w21;    //: /sn:0 {0}(710,270)(710,274){1}
//: {2}(712,276)(1064,276)(1064,-235)(98,-235)(98,646){3}
//: {4}(96,648)(74,648)(74,648)(61,648){5}
//: {6}(98,650)(98,749)(-449,749)(-449,793){7}
//: {8}(-447,795)(-437,795){9}
//: {10}(-451,795)(-459,795){11}
//: {12}(708,276)(705,276)(705,274)(700,274){13}
//: {14}(698,272)(698,264){15}
//: {16}(696,274)(686,274)(686,271){17}
//: {18}(686,267)(686,258){19}
//: {20}(684,269)(674,269)(674,266){21}
//: {22}(674,262)(674,253)(674,253)(674,252){23}
//: {24}(672,264)(662,264)(662,259){25}
//: {26}(662,255)(662,246){27}
//: {28}(660,257)(650,257)(650,251){29}
//: {30}(650,247)(650,240){31}
//: {32}(648,249)(638,249)(638,234){33}
wire w76;    //: /sn:0 {0}(941,2091)(931,2091){1}
//: {2}(929,2089)(929,2033)(1339,2033)(1339,1186){3}
//: {4}(1339,1182)(1339,587)(244,587)(244,270)(327,270)(327,274){5}
//: {6}(1337,1184)(1197,1184){7}
//: {8}(927,2091)(918,2091){9}
wire w374;    //: /sn:0 {0}(-377,1365)(-384,1365){1}
wire w340;    //: /sn:0 {0}(-165,1492)(-166,1492){1}
//: {2}(-168,1490)(-168,1430)(353,1430)(353,1158){3}
//: {4}(355,1156)(431,1156)(431,1156)(547,1156){5}
//: {6}(353,1154)(353,649)(155,649)(155,308)(355,308){7}
//: {8}(357,306)(357,304)(367,304){9}
//: {10}(369,306)(369,311)(369,311)(369,313){11}
//: {12}(369,302)(369,299)(379,299){13}
//: {14}(381,301)(381,304)(381,304)(381,307){15}
//: {16}(381,297)(381,294)(391,294){17}
//: {18}(393,296)(393,300)(393,300)(393,301){19}
//: {20}(393,292)(393,287)(403,287){21}
//: {22}(405,289)(405,295){23}
//: {24}(405,285)(405,280)(415,280){25}
//: {26}(417,282)(417,287)(417,287)(417,289){27}
//: {28}(417,278)(417,275)(427,275){29}
//: {30}(429,277)(429,280)(429,280)(429,283){31}
//: {32}(429,273)(429,270)(439,270){33}
//: {34}(441,272)(441,276)(441,276)(441,277){35}
//: {36}(441,268)(441,263)(451,263){37}
//: {38}(453,265)(453,270)(453,270)(453,271){39}
//: {40}(453,261)(453,258)(463,258){41}
//: {42}(465,260)(465,265){43}
//: {44}(465,256)(465,252)(477,252)(477,259){45}
//: {46}(357,310)(357,319){47}
//: {48}(-170,1492)(-187,1492){49}
wire w170;    //: /sn:0 {0}(863,1819)(856,1819){1}
wire w100;    //: /sn:0 {0}(1138,2239)(1128,2239){1}
//: {2}(1126,2237)(1126,2206)(1372,2206)(1372,1337){3}
//: {4}(1372,1333)(1372,552)(223,552)(223,-174)(534,-174)(534,-69)(529,-69){5}
//: {6}(1370,1335)(1348,1335)(1348,1334)(1197,1334){7}
//: {8}(1124,2239)(1116,2239){9}
wire w31;    //: /sn:0 {0}(1203,1658)(1194,1658){1}
//: {2}(1192,1656)(1192,1545)(1264,1545)(1264,866){3}
//: {4}(1264,862)(1264,669)(1001,669)(1001,95)(857,95)(857,80){5}
//: {6}(1262,864)(1197,864){7}
//: {8}(1190,1658)(1182,1658){9}
wire w24;    //: /sn:0 {0}(1010,1655)(995,1655){1}
//: {2}(993,1653)(993,1535)(1258,1535)(1258,836){3}
//: {4}(1258,832)(1258,675)(1007,675)(1007,-23)(802,-23){5}
//: {6}(1256,834)(1197,834){7}
//: {8}(991,1655)(984,1655){9}
wire w358;    //: /sn:0 {0}(-376,1075)(-383,1075){1}
wire w251;    //: /sn:0 {0}(925,2114)(918,2114){1}
wire w260;    //: /sn:0 {0}(600,2254)(593,2254){1}
wire w328;    //: /sn:0 {0}(-247,1220)(-252,1220){1}
wire w235;    //: /sn:0 {0}(601,2109)(594,2109){1}
wire w334;    //: /sn:0 {0}(-442,1217)(-447,1217){1}
wire w196;    //: /sn:0 {0}(97,1349)(89,1349){1}
//: {2}(87,1347)(87,1298)(333,1298)(333,1078){3}
//: {4}(335,1076)(421,1076)(421,1076)(547,1076){5}
//: {6}(333,1074)(333,661)(537,661)(537,470){7}
//: {8}(539,468)(545,468)(545,468)(541,468){9}
//: {10}(537,466)(537,462)(540,462)(540,458){11}
//: {12}(542,456)(548,456)(548,456)(544,456){13}
//: {14}(540,454)(540,449)(542,449)(542,445){15}
//: {16}(544,443)(550,443)(550,443)(546,443){17}
//: {18}(542,441)(542,436)(544,436)(544,432){19}
//: {20}(546,430)(553,430)(553,430)(549,430){21}
//: {22}(544,428)(544,419)(547,419)(547,419){23}
//: {24}(549,417)(556,417)(556,417)(552,417){25}
//: {26}(547,415)(547,411)(549,411)(549,406){27}
//: {28}(551,404)(558,404)(558,404)(554,404){29}
//: {30}(549,402)(549,397)(551,397)(551,393){31}
//: {32}(553,391)(560,391)(560,391)(556,391){33}
//: {34}(551,389)(551,385)(553,385)(553,381){35}
//: {36}(555,379)(562,379)(562,379)(558,379){37}
//: {38}(553,377)(553,373)(556,373)(556,369){39}
//: {40}(558,367)(565,367)(565,367)(561,367){41}
//: {42}(556,365)(556,360)(559,360)(559,356){43}
//: {44}(561,354)(568,354)(568,354)(564,354){45}
//: {46}(559,352)(559,341)(566,341){47}
//: {48}(85,1349)(73,1349){49}
wire w372;    //: /sn:0 {0}(143,1665)(138,1665){1}
wire w116;    //: /sn:0 {0}(397,1870)(444,1870){1}
//: {2}(446,1868)(446,1853)(446,1853)(446,1850){3}
//: {4}(448,1848)(477,1848){5}
//: {6}(481,1848)(527,1848)(527,1848)(539,1848){7}
//: {8}(543,1848)(604,1848){9}
//: {10}(608,1848)(615,1848)(615,1848)(671,1848){11}
//: {12}(675,1848)(707,1848)(707,1848)(738,1848){13}
//: {14}(742,1848)(788,1848)(788,1848)(800,1848){15}
//: {16}(804,1848)(865,1848){17}
//: {18}(869,1848)(919,1848)(919,1848)(930,1848){19}
//: {20}(934,1848)(941,1848)(941,1848)(997,1848){21}
//: {22}(1001,1848)(1033,1848)(1033,1848)(1064,1848){23}
//: {24}(1068,1848)(1114,1848)(1114,1848)(1126,1848){25}
//: {26}(1130,1848)(1160,1848)(1160,1848)(1194,1848)(1194,1825)(1203,1825){27}
//: {28}(1128,1846)(1128,1824)(1140,1824){29}
//: {30}(1066,1846)(1066,1823)(1076,1823){31}
//: {32}(999,1846)(999,1822)(1010,1822){33}
//: {34}(932,1846)(932,1821)(942,1821){35}
//: {36}(867,1846)(867,1820)(877,1820){37}
//: {38}(802,1846)(802,1819)(814,1819){39}
//: {40}(740,1846)(740,1818)(750,1818){41}
//: {42}(673,1846)(673,1817)(684,1817){43}
//: {44}(606,1846)(606,1816)(616,1816){45}
//: {46}(541,1846)(541,1815)(553,1815){47}
//: {48}(479,1846)(479,1814)(489,1814){49}
//: {50}(446,1846)(446,1705)(477,1705){51}
//: {52}(481,1705)(539,1705){53}
//: {54}(543,1705)(604,1705){55}
//: {56}(608,1705)(615,1705)(615,1705)(671,1705){57}
//: {58}(675,1705)(707,1705)(707,1705)(738,1705){59}
//: {60}(742,1705)(788,1705)(788,1705)(800,1705){61}
//: {62}(804,1705)(865,1705){63}
//: {64}(869,1705)(919,1705)(919,1705)(930,1705){65}
//: {66}(934,1705)(941,1705)(941,1705)(997,1705){67}
//: {68}(1001,1705)(1033,1705)(1033,1705)(1064,1705){69}
//: {70}(1068,1705)(1114,1705)(1114,1705)(1126,1705){71}
//: {72}(1130,1705)(1160,1705)(1160,1705)(1194,1705)(1194,1682)(1203,1682){73}
//: {74}(1128,1703)(1128,1681)(1140,1681){75}
//: {76}(1066,1703)(1066,1680)(1076,1680){77}
//: {78}(999,1703)(999,1679)(1010,1679){79}
//: {80}(932,1703)(932,1678)(942,1678){81}
//: {82}(867,1703)(867,1677)(877,1677){83}
//: {84}(802,1703)(802,1676)(814,1676){85}
//: {86}(740,1703)(740,1675)(750,1675){87}
//: {88}(673,1703)(673,1674)(684,1674){89}
//: {90}(606,1703)(606,1673)(616,1673){91}
//: {92}(541,1703)(541,1672)(553,1672){93}
//: {94}(479,1703)(479,1671)(489,1671){95}
//: {96}(446,1872)(446,1926)(446,1926)(446,1993){97}
//: {98}(448,1995)(476,1995){99}
//: {100}(480,1995)(526,1995)(526,1995)(538,1995){101}
//: {102}(542,1995)(603,1995){103}
//: {104}(607,1995)(614,1995)(614,1995)(670,1995){105}
//: {106}(674,1995)(706,1995)(706,1995)(737,1995){107}
//: {108}(741,1995)(787,1995)(787,1995)(799,1995){109}
//: {110}(803,1995)(864,1995){111}
//: {112}(868,1995)(918,1995)(918,1995)(929,1995){113}
//: {114}(933,1995)(940,1995)(940,1995)(996,1995){115}
//: {116}(1000,1995)(1032,1995)(1032,1995)(1063,1995){117}
//: {118}(1067,1995)(1113,1995)(1113,1995)(1125,1995){119}
//: {120}(1129,1995)(1193,1995)(1193,1972)(1202,1972){121}
//: {122}(1127,1993)(1127,1971)(1139,1971){123}
//: {124}(1065,1993)(1065,1970)(1075,1970){125}
//: {126}(998,1993)(998,1969)(1009,1969){127}
//: {128}(931,1993)(931,1968)(941,1968){129}
//: {130}(866,1993)(866,1967)(876,1967){131}
//: {132}(801,1993)(801,1966)(813,1966){133}
//: {134}(739,1993)(739,1965)(749,1965){135}
//: {136}(672,1993)(672,1964)(683,1964){137}
//: {138}(605,1993)(605,1963)(615,1963){139}
//: {140}(540,1993)(540,1962)(552,1962){141}
//: {142}(478,1993)(478,1961)(488,1961){143}
//: {144}(446,1997)(446,2140){145}
//: {146}(448,2142)(476,2142){147}
//: {148}(480,2142)(526,2142)(526,2142)(538,2142){149}
//: {150}(542,2142)(603,2142){151}
//: {152}(607,2142)(614,2142)(614,2142)(670,2142){153}
//: {154}(674,2142)(706,2142)(706,2142)(737,2142){155}
//: {156}(741,2142)(787,2142)(787,2142)(799,2142){157}
//: {158}(803,2142)(864,2142){159}
//: {160}(868,2142)(918,2142)(918,2142)(929,2142){161}
//: {162}(933,2142)(940,2142)(940,2142)(996,2142){163}
//: {164}(1000,2142)(1032,2142)(1032,2142)(1063,2142){165}
//: {166}(1067,2142)(1113,2142)(1113,2142)(1125,2142){167}
//: {168}(1129,2142)(1159,2142)(1159,2142)(1191,2142){169}
//: {170}(1195,2142)(1266,2142){171}
//: {172}(1193,2140)(1193,2119)(1202,2119){173}
//: {174}(1127,2140)(1127,2118)(1139,2118){175}
//: {176}(1065,2140)(1065,2117)(1075,2117){177}
//: {178}(998,2140)(998,2116)(1009,2116){179}
//: {180}(931,2140)(931,2115)(941,2115){181}
//: {182}(866,2140)(866,2114)(876,2114){183}
//: {184}(801,2140)(801,2113)(813,2113){185}
//: {186}(739,2140)(739,2112)(749,2112){187}
//: {188}(672,2140)(672,2111)(683,2111){189}
//: {190}(605,2140)(605,2110)(615,2110){191}
//: {192}(540,2140)(540,2109)(552,2109){193}
//: {194}(478,2140)(478,2108)(488,2108){195}
//: {196}(446,2144)(446,2287)(475,2287){197}
//: {198}(479,2287)(525,2287)(525,2287)(537,2287){199}
//: {200}(541,2287)(602,2287){201}
//: {202}(606,2287)(613,2287)(613,2287)(669,2287){203}
//: {204}(673,2287)(705,2287)(705,2287)(736,2287){205}
//: {206}(740,2287)(786,2287)(786,2287)(798,2287){207}
//: {208}(802,2287)(863,2287){209}
//: {210}(867,2287)(917,2287)(917,2287)(928,2287){211}
//: {212}(932,2287)(939,2287)(939,2287)(995,2287){213}
//: {214}(999,2287)(1031,2287)(1031,2287)(1062,2287){215}
//: {216}(1066,2287)(1112,2287)(1112,2287)(1124,2287){217}
//: {218}(1128,2287)(1192,2287)(1192,2264)(1201,2264){219}
//: {220}(1126,2285)(1126,2263)(1138,2263){221}
//: {222}(1064,2285)(1064,2262)(1074,2262){223}
//: {224}(997,2285)(997,2261)(1008,2261){225}
//: {226}(930,2285)(930,2260)(940,2260){227}
//: {228}(865,2285)(865,2259)(875,2259){229}
//: {230}(800,2285)(800,2258)(812,2258){231}
//: {232}(738,2285)(738,2257)(748,2257){233}
//: {234}(671,2285)(671,2256)(682,2256){235}
//: {236}(604,2285)(604,2255)(614,2255){237}
//: {238}(539,2285)(539,2254)(551,2254){239}
//: {240}(477,2285)(477,2253)(487,2253){241}
wire w98;    //: /sn:0 {0}(926,1677)(919,1677){1}
wire w18;    //: /sn:0 {0}(397,1682)(281,1682)(281,1767){1}
wire w243;    //: /sn:0 {0}(664,2110)(657,2110){1}
wire w118;    //: /sn:0 {0}(10,825)(-6,825){1}
wire w212;    //: /sn:0 {0}(862,1966)(855,1966){1}
wire w68;    //: /sn:0 {0}(615,2086)(603,2086){1}
//: {2}(601,2084)(601,2008)(1329,2008)(1329,1136){3}
//: {4}(1329,1132)(1329,597)(254,597)(254,440)(390,440)(390,430)(400,430){5}
//: {6}(1327,1134)(1197,1134){7}
//: {8}(599,2086)(594,2086){9}
wire w371;    //: /sn:0 {0}(-182,1368)(-187,1368){1}
wire w59;    //: /sn:0 {0}(1009,1945)(1000,1945){1}
//: {2}(998,1943)(998,1889)(1314,1889)(1314,1076){3}
//: {4}(1314,1072)(1314,613)(553,613)(553,483)(563,483){5}
//: {6}(1312,1074)(1197,1074){7}
//: {8}(996,1945)(983,1945){9}
wire w123;    //: /sn:0 {0}(991,1678)(984,1678){1}
wire w62;    //: /sn:0 {0}(1139,1947)(1133,1947){1}
//: {2}(1131,1945)(1131,1897)(1318,1897)(1318,1096){3}
//: {4}(1318,1092)(1318,609)(501,609)(501,480)(511,480){5}
//: {6}(1316,1094)(1197,1094){7}
//: {8}(1129,1947)(1117,1947){9}
wire w85;    //: /sn:0 {0}(863,1676)(856,1676){1}
wire w185;    //: /sn:0 {0}(1057,1822)(1052,1822){1}
wire w11;    //: /sn:0 {0}(1118,1657)(1124,1657){1}
//: {2}(1128,1657)(1140,1657){3}
//: {4}(1126,1655)(1126,1542)(1262,1542)(1262,856){5}
//: {6}(1262,852)(1262,671)(1003,671)(1003,54)(891,54)(891,72)(845,72)(845,43){7}
//: {8}(1260,854)(1197,854){9}
wire w137;    //: /sn:0 {0}(-715,814)(-720,814){1}
wire w70;    //: /sn:0 {0}(657,2087)(670,2087){1}
//: {2}(674,2087)(683,2087){3}
//: {4}(672,2085)(672,2013)(1331,2013)(1331,1146){5}
//: {6}(1331,1142)(1331,595)(252,595)(252,387)(376,387)(376,397){7}
//: {8}(1329,1144)(1197,1144){9}
wire w193;    //: /sn:0 {0}(355,361)(355,351)(250,351)(250,593)(1333,593)(1333,1152){1}
//: {2}(1331,1154)(1197,1154){3}
//: {4}(1333,1156)(1333,2018)(735,2018)(735,2086){5}
//: {6}(737,2088)(749,2088){7}
//: {8}(733,2088)(725,2088){9}
wire w110;    //: /sn:0 {0}(1189,1681)(1182,1681){1}
wire w189;    //: /sn:0 {0}(536,1814)(531,1814){1}
wire w206;    //: /sn:0 {0}(796,1965)(791,1965){1}
wire w13;    //: /sn:0 {0}(1197,874)(1264,874){1}
//: {2}(1266,872)(1266,667)(999,667)(999,116)(866,116)(866,103){3}
//: {4}(1266,876)(1266,1549)(1259,1549)(1259,1657){5}
//: {6}(1257,1659)(1245,1659){7}
//: {8}(1259,1661)(1259,1710)(479,1710)(479,1790)(489,1790){9}
wire w353;    //: /sn:0 {0}(144,1373)(139,1373){1}
wire w88;    //: /sn:0 {0}(-388,819)(-395,819){1}
wire w5;    //: /sn:0 {0}(553,1648)(542,1648){1}
//: {2}(540,1646)(540,1593){3}
//: {4}(540,1589)(540,1504)(1244,1504)(1244,766){5}
//: {6}(1244,762)(1244,689)(1021,689)(1021,-189)(610,-189)(610,-72)(607,-72){7}
//: {8}(1242,764)(1197,764){9}
//: {10}(538,1591)(431,1591)(431,1740)(-634,1740)(-634,1098)(-604,1098){11}
//: {12}(538,1648)(531,1648){13}
wire w48;    //: /sn:0 {0}(1052,1799)(1065,1799){1}
//: {2}(1069,1799)(1076,1799){3}
//: {4}(1067,1797)(1067,1753)(1288,1753)(1288,966){5}
//: {6}(1288,962)(1288,641)(1041,641)(1041,353)(856,353)(856,341){7}
//: {8}(1286,964)(1197,964){9}
wire w47;    //: /sn:0 {0}(984,1798)(996,1798){1}
//: {2}(1000,1798)(1010,1798){3}
//: {4}(998,1796)(998,1749)(1286,1749)(1286,956){5}
//: {6}(1286,952)(1286,643)(1039,643)(1039,324)(865,324)(865,316){7}
//: {8}(1284,954)(1197,954){9}
wire w26;    //: /sn:0 {0}(-824,848)(-818,848)(-818,643)(-812,643){1}
wire w342;    //: /sn:0 {0}(79,1082)(74,1082){1}
//: enddecls

  //: joint g8 (w119) @(1259, 2228) /w:[ 2 4 -1 1 ]
  //: joint g1883 (w120) @(-113, 1638) /w:[ 10 9 12 -1 ]
  //: joint g1482 (w352) @(337, 140) /anc:1 /w:[ 3 -1 4 14 ]
  //: joint g1397 (w196) @(544, 430) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g611 (w265) @(395,61) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1783 (w108) @(212, 1643) /w:[ 46 45 48 -1 ]
  //: joint g2045 (w297) @(331, 1066) /w:[ 4 6 -1 3 ]
  //: joint g139 (w153) @(734, -25) /anc:1 /w:[ 11 -1 12 14 ]
  //: joint g659 (w202) @(450, 362) /anc:1 /w:[ 27 -1 28 30 ]
  //: joint g465 (w28) @(610, 5) /anc:1 /w:[ 29 30 32 -1 ]
  D_FF g1841 (.D(w113), .CP(w34), .Q(w35), .NQ(w371));   //: @(-228, 1331) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>135 Ro0<49 Ro1<1 ]
  //: joint g521 (w341) @(742, 55) /anc:1 /w:[ 31 -1 32 34 ]
  //: LED g529 (w341) @(749,33) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: joint g658 (w202) @(468, 340) /anc:1 /w:[ 35 -1 36 38 ]
  //: joint g813 (w0) @(419, 351) /anc:1 /w:[ 17 18 -1 20 ]
  //: LED g831 (w120) @(410,-10) /sn:0 /R:1 /anc:1 /w:[ 15 ] /type:0
  D_FF g1731 (.D(w0), .CP(w34), .Q(w204), .NQ(w285));   //: @(-294, 1477) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>189 Ro0<49 Ro1<1 ]
  //: LED g932 (w211) @(400,221) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g1366 (w116) @(801, 2142) /w:[ 158 184 157 -1 ]
  //: joint g720 (w298) @(703, 334) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g982 (w103) @(767, 149) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g1398 (w304) @(548,377) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g508 (w87) @(741, 22) /anc:1 /w:[ 19 -1 20 22 ]
  //: joint g1305 (w134) @(635, -33) /anc:1 /w:[ -1 15 16 18 ]
  //: joint g621 (w183) @(736, 427) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g1734 (w34) @(-438, 1398) /w:[ 102 140 101 -1 ]
  //: joint g2023 (w120) @(384, 1286) /w:[ 6 5 -1 8 ]
  //: joint g1089 (w283) @(414, 228) /anc:1 /w:[ 29 30 32 -1 ]
  //: joint g38 (w10) @(805, 1652) /w:[ 1 2 8 -1 ]
  //: LED g1544 (w163) @(643,-20) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g307 (w186) @(692,387) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g568 (w181) @(803,381) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g665 (w202) @(434,395) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g850 (w120) @(460, 32) /anc:1 /w:[ 25 26 -1 28 ]
  //: LED g393 (w22) @(626,255) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  _GGOR2 #(6) g1788 (.I0(w115), .I1(w112), .Z(w34));   //: @(-537,925) /sn:0 /w:[ 1 1 95 ]
  //: joint g1655 (w46) @(866, 1796) /w:[ 2 4 1 -1 ]
  //: joint g1592 (w174) @(771, 267) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g792 (w16) @(-319, 848) /w:[ 16 30 15 -1 ]
  //: joint g1706 (w121) @(-625, 1136) /w:[ -1 1 2 4 ]
  //: LED g969 (w64) @(581,-7) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  D_FF g885 (.D(w40), .CP(w116), .Q(w44), .NQ(w162));   //: @(751, 1781) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>41 Ro0<0 Ro1<1 ]
  //: joint g1530 (w163) @(640, 56) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1059 (w111) @(862, 165) /anc:1 /w:[ -1 4 6 3 ]
  //: joint g2034 (w356) @(357, 1176) /w:[ 4 6 -1 3 ]
  //: joint g1917 (w15) @(1254, 814) /w:[ -1 4 6 3 ]
  //: LED g1498 (w357) @(696,-35) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g902 (w89) @(826, 194) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g917 (w33) @(620,442) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1690 (w86) @(602, 2231) /w:[ 1 2 8 -1 ]
  //: joint g1508 (w151) @(679, -31) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g696 (w332) @(764, 107) /anc:1 /w:[ 31 32 -1 34 ]
  //: LED g732 (w204) @(437,312) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g818 (w0) @(495,297) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g834 (w120) @(479, 53) /anc:1 /w:[ 33 34 -1 36 ]
  //: joint g886 (w16) @(-511, 848) /w:[ 10 36 9 -1 ]
  //: LED g93 (w100) @(522,-69) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: LED g852 (w111) @(761,173) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g768 (w296) @(517, 63) /anc:1 /w:[ 39 40 -1 42 ]
  //: LED g26 (w19) @(688,204) /sn:0 /anc:1 /w:[ 17 ] /type:0
  D_FF g1372 (.D(w75), .CP(w116), .Q(w74), .NQ(w237));   //: @(814, 2076) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>185 Ro0<9 Ro1<1 ]
  //: LED g1546 (w163) @(626,69) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: LED g1395 (w304) @(542,402) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1257 (w297) @(564, 443) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1206 (w141) @(543, -30) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g1679 (w50) @(1130, 1800) /w:[ 2 4 1 -1 ]
  //: LED g34 (w20) @(600,143) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g963 (w64) @(584,30) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g1759 (w352) @(280, 1499) /w:[ -1 9 10 12 ]
  //: comment g1989 @(325,320)
  //: /line:"<h1 color=blue>8</h1>"
  //: /end
  //: joint g1242 (w171) @(837, 239) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g267 (w317) @(465, 436) /anc:1 /w:[ 11 -1 12 14 ]
  //: joint g1878 (w28) @(-438, 1051) /w:[ 1 2 52 -1 ]
  //: joint g1115 (w108) @(563, -46) /anc:1 /w:[ 7 8 10 -1 ]
  //: joint g523 (w341) @(751, 44) /anc:1 /w:[ 27 -1 28 30 ]
  //: LED g1120 (w108) @(572,56) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1695 (w116) @(446, 1995) /w:[ 98 97 -1 144 ]
  //: joint g1480 (w219) @(339, 116) /anc:1 /w:[ 10 -1 9 48 ]
  //: joint g451 (w28) @(610, -46) /anc:1 /w:[ 13 14 16 -1 ]
  //: LED g325 (w186) @(710,423) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: LED g397 (w22) @(632,267) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1359 (w116) @(739, 1995) /w:[ 108 134 107 -1 ]
  D_FF g1616 (.D(w68), .CP(w116), .Q(w70), .NQ(w243));   //: @(616, 2073) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>191 Ro0<0 Ro1<1 ]
  //: joint g1036 (w360) @(515, -38) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g577 (w287) @(746, 321) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g1284 (w215) @(375,181) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: joint g433 (w19) @(725, 221) /anc:1 /w:[ 3 4 6 -1 ]
  //: joint g280 (w317) @(476, 412) /anc:1 /w:[ 19 -1 20 22 ]
  //: joint g1220 (w116) @(999, 1848) /w:[ 22 32 21 -1 ]
  //: joint g1791 (w34) @(-306, 1545) /w:[ 154 188 153 -1 ]
  //: joint g1873 (w34) @(-372, 1251) /w:[ 33 34 36 -1 ]
  //: joint g1013 (w207) @(408, 267) /anc:1 /w:[ 21 22 24 -1 ]
  //: LED g752 (w296) @(491,39) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g1056 (w111) @(824, 171) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g663 (w202) @(470,351) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g1302 (w215) @(401,183) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g2039 (w202) @(347, 1126) /w:[ 4 6 -1 3 ]
  //: joint g469 (w28) @(610, -33) /anc:1 /w:[ 17 18 20 -1 ]
  //: LED g1118 (w108) @(553,-46) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g717 (w298) @(712, 345) /anc:1 /w:[ 35 36 -1 38 ]
  //: joint g1524 (w163) @(657, -33) /anc:1 /w:[ -1 15 16 18 ]
  //: joint g1667 (w55) @(737, 1941) /w:[ 1 2 8 -1 ]
  //: LED g1196 (w141) @(552,33) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: LED g1249 (w171) @(850,228) /sn:0 /anc:1 /w:[ 13 ] /type:0
  D_FF g1343 (.D(w58), .CP(w116), .Q(w59), .NQ(w200));   //: @(942, 1931) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>129 Ro0<9 Ro1<1 ]
  //: joint g1919 (w6) @(1248, 784) /w:[ -1 4 6 3 ]
  //: joint g2050 (w314) @(321, 1016) /w:[ 4 6 -1 3 ]
  //: LED g95 (w119) @(575,-72) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  D_FF g1815 (.D(w177), .CP(w34), .Q(w286), .NQ(w362));   //: @(33, 1188) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>11 Ro0<49 Ro1<1 ]
  //: joint g1934 (w48) @(1288, 964) /w:[ -1 6 8 5 ]
  //: LED g24 (w22) @(656,315) /sn:0 /R:3 /anc:1 /w:[ 0 ] /type:0
  //: joint g1687 (w91) @(865, 2235) /w:[ 2 4 1 -1 ]
  //: joint g1743 (w196) @(87, 1349) /w:[ 1 2 48 -1 ]
  D_FF g1223 (.D(w109), .CP(w16), .Q(w20), .NQ(w137));   //: @(-761, 777) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>45 Ro0<0 Ro1<1 ]
  //: joint g594 (w183) @(719, 404) /anc:1 /w:[ 19 20 -1 22 ]
  //: LED g251 (w29) @(512,202) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g204 (w169) @(839, 216) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g303 (w286) @(734, 293) /anc:1 /w:[ -1 44 46 43 ]
  //: joint g332 (w186) @(676, 387) /anc:1 /w:[ 27 28 -1 30 ]
  //: joint g1503 (w163) @(648, 19) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g431 (w22) @(634, 315) /anc:1 /w:[ 1 2 -1 24 ]
  //: joint g97 (w153) @(688, 71) /anc:1 /w:[ 43 -1 44 46 ]
  //: LED g895 (w89) @(826,184) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g239 (w224) @(408,104) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1536 (w151) @(642,58) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g970 (w64) @(578,-46) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g896 (w89) @(751, 200) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g1114 (w108) @(558,-20) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g1209 (w174) @(759,250) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g936 (w211) @(450, 207) /anc:1 /w:[ 41 42 44 -1 ]
  //: joint g1816 (w356) @(-49, 1494) /w:[ 1 2 48 -1 ]
  //: comment g1986 @(726,466)
  //: /line:"<h1 color=blue>5</h1>"
  //: /end
  //: LED g1571 (w174) @(796,261) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: SWITCH g1979 (w117) @(343,-73) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:0
  //: joint g709 (w332) @(799, 85) /anc:1 /w:[ 19 20 -1 22 ]
  //: joint g1214 (w174) @(848, 286) /anc:1 /w:[ 7 8 10 -1 ]
  //: LED g319 (w25) @(565,268) /sn:0 /R:3 /anc:1 /w:[ 23 ] /type:0
  //: joint g991 (w314) @(643, 347) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g561 (w201) @(444,432) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1639 (w116) @(1126, 2287) /w:[ 218 220 217 -1 ]
  //: joint g960 (w64) @(589, -33) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g206 (w274) @(463,202) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g274 (w317) @(529,340) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g294 (w286) @(758, 304) /anc:1 /w:[ 35 -1 36 38 ]
  D_FF g1607 (.D(w70), .CP(w116), .Q(w193), .NQ(w239));   //: @(684, 2074) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>189 Ro0<9 Ro1<1 ]
  //: joint g1447 (w352) @(426, 156) /anc:1 /w:[ 37 38 40 -1 ]
  //: joint g472 (w300) @(589, 456) /anc:1 /w:[ 7 8 10 -1 ]
  //: joint g871 (w116) @(999, 1705) /w:[ 68 78 67 -1 ]
  //: LED g1098 (w283) @(350,250) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: joint g1256 (w297) @(568, 404) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1182 (w356) @(392,262) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g904 (w89) @(788,187) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g842 (w120) @(432, 0) /anc:1 /w:[ 2 1 -1 16 ]
  //: joint g1104 (w283) @(389, 232) /anc:1 /w:[ 21 22 24 -1 ]
  //: joint g1956 (w76) @(1339, 1184) /w:[ -1 4 6 3 ]
  //: LED g493 (w87) @(680,90) /sn:0 /R:1 /anc:1 /w:[ 43 ] /type:0
  //: LED g864 (w360) @(541,49) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1727 (w34) @(148, 1690) /w:[ 218 220 217 -1 ]
  //: joint g815 (w0) @(408, 362) /anc:1 /w:[ 13 14 -1 16 ]
  //: LED g758 (w296) @(483,27) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g685 (w228) @(408,36) /sn:0 /R:2 /anc:1 /w:[ 17 ] /type:0
  //: LED g276 (w317) @(523,352) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g340 (w186) @(722,447) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  D_FF g1338 (.D(w13), .CP(w116), .Q(w132), .NQ(w189));   //: @(490, 1777) /sz:(40, 56) /sn:0 /p:[ Li0>9 Li1>49 Ro0<9 Ro1<1 ]
  //: joint g1630 (w116) @(671, 2287) /w:[ 204 234 203 -1 ]
  //: SWITCH g798 (w104) @(254,-73) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:0
  //: joint g629 (w183) @(728, 416) /anc:1 /w:[ 15 16 -1 18 ]
  //: joint g567 (w181) @(748, 347) /anc:1 /w:[ 31 -1 32 34 ]
  //: joint g1112 (w108) @(573, 5) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g482 (w300) @(589, 417) /anc:1 /w:[ 19 20 22 -1 ]
  D_FF g797 (.D(w23), .CP(w116), .Q(w5), .NQ(w43));   //: @(490, 1634) /sz:(40, 56) /sn:0 /p:[ Li0>1 Li1>95 Ro0<13 Ro1<1 ]
  //: LED g202 (w274) @(362,202) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g446 (w340) @(417, 280) /anc:1 /w:[ 25 26 -1 28 ]
  //: LED g1295 (w215) @(414,184) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g94 (w96) @(547,-72) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: joint g899 (w89) @(788, 197) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g287 (w286) @(842, 345) /anc:1 /w:[ 7 8 10 -1 ]
  D_FF g1360 (.D(w60), .CP(w116), .Q(w62), .NQ(w220));   //: @(1076, 1933) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>125 Ro0<9 Ro1<1 ]
  //: joint g1010 (w207) @(421, 262) /anc:1 /w:[ 25 26 28 -1 ]
  //: LED g458 (w28) @(600,55) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g1940 (w56) @(1304, 1024) /w:[ -1 4 6 3 ]
  D_FF g800 (.D(w5), .CP(w116), .Q(w3), .NQ(w102));   //: @(554, 1635) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>93 Ro0<9 Ro1<1 ]
  //: LED g345 (w67) @(504,151) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: LED g1464 (w290) @(458,145) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  //: joint g91 (w116) @(541, 1705) /w:[ 54 92 53 -1 ]
  D_FF g1370 (.D(w66), .CP(w116), .Q(w68), .NQ(w235));   //: @(553, 2072) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>193 Ro0<9 Ro1<1 ]
  //: LED g269 (w317) @(535,328) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: joint g639 (w181) @(759, 356) /anc:1 /w:[ 27 -1 28 30 ]
  //: LED g952 (w64) @(582,5) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: joint g1945 (w59) @(1314, 1074) /w:[ -1 4 6 3 ]
  //: joint g1623 (w65) @(1258, 1949) /w:[ -1 2 1 8 ]
  //: joint g1699 (w141) @(148, 1642) /w:[ 46 45 48 -1 ]
  _GGAND2 #(6) g1866 (.I0(w117), .I1(w121), .Z(w116));   //: @(387,1870) /sn:0 /w:[ 1 7 0 ]
  //: joint g1259 (w297) @(573, 354) /anc:1 /w:[ 43 44 46 -1 ]
  //: LED g213 (w274) @(450,202) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  D_FF g889 (.D(w21), .CP(w16), .Q(w22), .NQ(w88));   //: @(-436, 782) /sz:(40, 56) /sn:0 /p:[ Li0>9 Li1>35 Ro0<33 Ro1<1 ]
  //: LED g1047 (w360) @(526,12) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g203 (w41) @(599,304) /sn:0 /R:3 /anc:1 /w:[ 15 ] /type:0
  D_FF g803 (.D(w15), .CP(w116), .Q(w14), .NQ(w98));   //: @(878, 1640) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>83 Ro0<9 Ro1<1 ]
  //: joint g1293 (w215) @(414, 172) /anc:1 /w:[ 29 30 32 -1 ]
  //: LED g1271 (w297) @(581,391) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g511 (w87) @(732, 34) /anc:1 /w:[ 23 -1 24 26 ]
  //: LED g1557 (w177) @(827,295) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g1160 (w113) @(637, 376) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g855 (w113) @(644,364) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: LED g847 (w120) @(420,0) /sn:0 /R:1 /anc:1 /w:[ 0 ] /type:0
  D_FF g1362 (.D(w59), .CP(w116), .Q(w60), .NQ(w223));   //: @(1010, 1932) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>127 Ro0<9 Ro1<1 ]
  //: joint g1668 (w56) @(672, 1940) /w:[ 1 2 8 -1 ]
  //: joint g1918 (w24) @(1258, 834) /w:[ -1 4 6 3 ]
  //: joint g1528 (w163) @(643, 43) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g1429 (w196) @(563,391) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g1026 (w207) @(471,252) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  //: LED g57 (w56) @(705,472) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g1506 (w163) @(646, 31) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1282 (w215) @(375, 169) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g484 (w300) @(589, 380) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1971 (w100) @(1372, 1335) /w:[ -1 4 6 3 ]
  //: joint g2074 (w163) @(263, 776) /w:[ 4 6 -1 3 ]
  //: joint g849 (w120) @(507, 86) /anc:1 /w:[ 45 46 -1 48 ]
  //: LED g1049 (w360) @(531,25) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: LED g1111 (w108) @(555,-33) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g674 (w228) @(452, 61) /anc:1 /w:[ 31 -1 32 34 ]
  //: LED g535 (w183) @(710,369) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g839 (w120) @(498, 75) /anc:1 /w:[ 41 42 -1 44 ]
  //: joint g1471 (w352) @(451, 162) /anc:1 /w:[ 45 46 48 -1 ]
  //: joint g1244 (w171) @(785, 234) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1116 (w108) @(568, -20) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g181 (w169) @(801, 216) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1535 (w151) @(663, 33) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g215 (w274) @(413,202) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  _GGOR2 #(6) g1640 (.I0(w7), .I1(w64), .Z(w2));   //: @(-653,1180) /sn:0 /R:1 /w:[ 9 49 0 ]
  //: joint g1710 (w21) @(-449, 795) /w:[ 8 7 10 -1 ]
  //: LED g827 (w0) @(398,383) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g1492 (w151) @(676,-56) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  D_FF g1739 (.D(w163), .CP(w34), .Q(w151), .NQ(w294));   //: @(-293, 1040) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>87 Ro0<49 Ro1<1 ]
  //: joint g1741 (w34) @(-177, 1398) /w:[ 110 132 109 -1 ]
  //: joint g1744 (w357) @(-173, 1055) /w:[ 1 2 48 -1 ]
  D_FF g1831 (.D(w202), .CP(w34), .Q(w0), .NQ(w367));   //: @(-362, 1476) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>191 Ro0<49 Ro1<1 ]
  _GGMUX2 #(40, 40) g1693 (.I0(w121), .I1(w30), .S(fdbk60), .Z(w26));   //: @(-837,848) /sn:0 /R:1 /delay:" 40 40" /w:[ 3 0 5 0 ] /ss:0 /do:0
  //: LED g541 (w228) @(386,18) /sn:0 /R:2 /anc:1 /w:[ 49 ] /type:0
  //: LED g30 (w13) @(866,96) /sn:0 /anc:1 /w:[ 3 ] /type:0
  //: LED g323 (w25) @(547,304) /sn:0 /R:3 /anc:1 /w:[ 11 ] /type:0
  //: joint g817 (w0) @(440, 333) /anc:1 /w:[ 25 26 -1 28 ]
  //: joint g1685 (w97) @(1063, 2238) /w:[ 1 2 8 -1 ]
  //: joint g2028 (w219) @(374, 1236) /w:[ 6 8 -1 5 ]
  //: LED g1439 (w290) @(360,106) /sn:0 /R:2 /anc:1 /w:[ 13 ] /type:0
  //: joint g514 (w87) @(701, 81) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g1138 (w330) @(859, 140) /anc:1 /w:[ -1 8 10 7 ]
  //: joint g771 (w296) @(457, -30) /anc:1 /w:[ 10 9 48 -1 ]
  D_FF g1231 (.D(w41), .CP(w16), .Q(w25), .NQ(w146));   //: @(-308, 784) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>31 Ro0<33 Ro1<1 ]
  //: LED g37 (w156) @(878,180) /sn:0 /anc:1 /w:[ 3 ] /type:0
  //: LED g1553 (w173) @(748,232) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1155 (w113) @(652, 426) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g1130 (w330) @(834,136) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g374 (w340) @(405,302) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g428 (w32) @(575, 128) /anc:1 /w:[ 15 16 -1 18 ]
  //: joint g1642 (w116) @(865, 2287) /w:[ 210 228 209 -1 ]
  //: joint g1904 (w41) @(102, 628) /w:[ -1 4 30 3 ]
  //: joint g1821 (w87) @(-50, 1057) /w:[ 46 45 48 -1 ]
  //: joint g218 (w274) @(437, 192) /anc:1 /w:[ 38 -1 37 44 ]
  //: joint g314 (w25) @(530, 304) /anc:1 /w:[ 10 12 9 -1 ]
  //: joint g1394 (w304) @(533, 389) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1949 (w65) @(1322, 1114) /w:[ -1 4 6 3 ]
  //: LED g766 (w296) @(444,-30) /sn:0 /R:1 /anc:1 /w:[ 49 ] /type:0
  //: LED g50 (w50) @(843,370) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g1086 (w35) @(636,404) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g1038 (w360) @(536,37) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g266 (w317) @(459, 448) /anc:1 /w:[ 8 10 -1 7 ]
  //: LED g19 (w10) @(707,-61) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: joint g638 (w181) @(737, 338) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g1514 (w151) @(657,8) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: joint g736 (w204) @(414, 312) /anc:1 /w:[ 21 22 -1 24 ]
  //: joint g1538 (w357) @(709, -47) /anc:1 /w:[ 8 7 -1 10 ]
  D_FF g1233 (.D(w73), .CP(w116), .Q(w47), .NQ(w157));   //: @(943, 1784) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>35 Ro0<0 Ro1<1 ]
  //: LED g984 (w103) @(804,124) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1807 (w134) @(-374, 1052) /w:[ 1 2 48 -1 ]
  //: LED g1247 (w171) @(811,224) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g724 (w298) @(733,356) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g837 (w120) @(470, 42) /anc:1 /w:[ 29 30 -1 32 ]
  //: joint g1736 (w177) @(20, 1201) /w:[ 1 2 48 -1 ]
  //: joint g1779 (w34) @(-373, 1545) /w:[ 152 190 151 -1 ]
  //: LED g524 (w341) @(713,77) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g865 (w64) @(592, 5) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g616 (w265) @(383,53) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: joint g2053 (w298) @(311, 986) /w:[ 4 6 -1 3 ]
  //: LED g1515 (w357) @(667,39) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g1444 (w352) @(414, 154) /anc:1 /w:[ 33 34 36 -1 ]
  //: joint g231 (w41) @(586, 304) /anc:1 /w:[ 14 16 -1 13 ]
  //: joint g2036 (w340) @(353, 1156) /w:[ 4 6 -1 3 ]
  //: joint g221 (w41) @(586, 317) /anc:1 /w:[ 10 12 -1 9 ]
  //: joint g2018 (w108) @(394, 1336) /w:[ 1 2 -1 44 ]
  //: joint g1493 (w151) @(654, 58) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1443 (w290) @(434, 123) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g1164 (w113) @(636,338) /sn:0 /R:3 /anc:1 /w:[ 43 ] /type:0
  //: joint g866 (w111) @(786, 178) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g755 (w296) @(510, 51) /anc:1 /w:[ 35 36 -1 38 ]
  //: LED g1066 (w111) @(799,166) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g249 (w29) @(550,202) /sn:0 /R:2 /anc:1 /w:[ 17 ] /type:0
  //: joint g1881 (w34) @(-111, 1108) /w:[ 62 80 61 -1 ]
  //: joint g0 (w7) @(54, 1872) /w:[ 1 2 8 -1 ]
  //: comment Welcome @(-452,314)
  //: /line:"<h1 color=Yellow3>Welcome to LEDClock </h1>"
  //: /line:"<font size=6 color=\"firebrick\">Computer Architecture </font>"
  //: /line:"<font size=6 color=\"firebrick\">Prof. Alessandro Bogliolo</font>"
  //: /line:""
  //: /line:"<font size=6 color=\"firebrick\">Individual Project</font>"
  //: /line:"<font size=4 color=\"firebrick\">Student Pirazzi Fulvio</font>"
  //: /line:"<font size=4 color=\"firebrick\">Serial numbers # 266093</font>"
  //: /line:"<font size=4 color=\"firebrick\">Year of enrolment second</font>"
  //: /line:""
  //: /line:"<font size=4 color=black>LEDClock provides a digital and analog clocks.</font>"
  //: /line:"<font size=4 color=black>In the frame Digital clock are 3 bottons:</font>"
  //: /line:"<font size=4 color=black>use [+1 h] and [+1 m] in order to increase the time</font>"
  //: /line:"<font size=4 color=black> [Run] to stop-continue</font>"
  //: /end
  //: LED g1376 (w304) @(560,339) /sn:0 /R:3 /anc:1 /w:[ 43 ] /type:0
  //: joint g919 (w33) @(606, 391) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1299 (w215) @(388, 170) /anc:1 /w:[ 21 22 24 -1 ]
  //: LED g1245 (w171) @(798,223) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g1579 (w177) @(777, 287) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1092 (w283) @(401, 230) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g395 (w22) @(617, 267) /anc:1 /w:[ 16 -1 18 15 ]
  //: comment g1978 @(868,49)
  //: /line:"<h1 color=blue>2</h1>"
  //: /end
  //: joint g1031 (w360) @(556, 62) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g86 (w19) @(725,204) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: LED g1436 (w219) @(466,163) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g346 (w233) @(501,8) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g655 (w202) @(425,406) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g59 (w69) @(650,481) /sn:0 /R:3 /anc:1 /w:[ 0 ] /type:0
  //: LED g1310 (w151) @(654,21) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g1488 (w290) @(397, 110) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g576 (w287) @(794, 353) /anc:1 /w:[ 19 -1 20 22 ]
  //: LED g592 (w287) @(818,355) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g1198 (w141) @(537, -55) /anc:1 /w:[ -1 3 4 6 ]
  //: LED g122 (w160) @(832,87) /sn:0 /anc:1 /w:[ 13 ] /type:0
  D_FF g1802 (.D(w340), .CP(w34), .Q(w207), .NQ(w355));   //: @(-164, 1479) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>185 Ro0<49 Ro1<1 ]
  //: LED g670 (w202) @(506,308) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  D_FF g794 (.D(w9), .CP(w116), .Q(w10), .NQ(w39));   //: @(751, 1638) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>87 Ro0<9 Ro1<1 ]
  //: LED g244 (w224) @(468,133) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: joint g1660 (w64) @(278, 1644) /w:[ -1 2 1 48 ]
  //: LED g119 (w153) @(670,71) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g921 (w33) @(612,341) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g15 (w149) @(622,167) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: joint g578 (w287) @(770, 337) /anc:1 /w:[ 27 -1 28 30 ]
  //: joint g1573 (w173) @(824, 259) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g1513 (w151) @(666, 21) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g923 (w33) @(615,379) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g757 (w296) @(465, -19) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g857 (w89) @(801, 196) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g2040 (w201) @(345, 1116) /w:[ 4 6 -1 3 ]
  //: LED g1279 (w196) @(548,468) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: LED g1080 (w35) @(627,353) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: LED g390 (w166) @(640,183) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g88 (w90) @(434,-42) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  //: joint g499 (w116) @(673, 1705) /w:[ 58 88 57 -1 ]
  //: joint g1797 (w35) @(-178, 1345) /w:[ 1 2 48 -1 ]
  //: joint g1809 (w34) @(-437, 1108) /w:[ 52 90 51 -1 ]
  //: joint g1537 (w151) @(672, -5) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g597 (w265) @(419, 62) /anc:1 /w:[ 21 -1 22 24 ]
  //: joint g607 (w265) @(467, 95) /anc:1 /w:[ 37 -1 38 40 ]
  //: joint g763 (w296) @(526, 75) /anc:1 /w:[ 43 44 -1 46 ]
  //: joint g369 (w233) @(509, -4) /anc:1 /w:[ 19 20 -1 22 ]
  //: LED g285 (w317) @(476,448) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g5 (w5) @(540, 1648) /w:[ 1 2 12 -1 ]
  //: joint g1855 (w304) @(153, 1350) /w:[ 46 45 48 -1 ]
  //: joint g2071 (w153) @(269, 806) /w:[ 4 6 -1 3 ]
  //: LED g1187 (w356) @(416,255) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: joint g1419 (w71) @(490, 457) /anc:1 /w:[ 8 10 -1 7 ]
  //: joint g1892 (w330) @(-435, 1194) /w:[ 1 2 48 -1 ]
  //: LED g626 (w183) @(734,404) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g1470 (w290) @(410, 114) /anc:1 /w:[ 23 24 26 -1 ]
  D_FF g1612 (.D(w79), .CP(w116), .Q(w77), .NQ(w242));   //: @(1140, 2081) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>175 Ro0<0 Ro1<1 ]
  //: joint g1875 (w34) @(-500, 1398) /w:[ 100 142 99 -1 ]
  //: joint g956 (w64) @(596, 55) /anc:1 /w:[ 43 44 46 -1 ]
  //: LED g779 (w339) @(794,33) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g1574 (w174) @(771,255) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: LED g18 (w9) @(680,-70) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  //: LED g739 (w204) @(390,343) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: LED g191 (w169) @(801,204) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g1156 (w113) @(647,376) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g1523 (w357) @(657,63) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: joint g336 (w67) @(504, 134) /anc:1 /w:[ 8 7 -1 26 ]
  //: joint g1333 (w116) @(740, 1848) /w:[ 14 40 13 -1 ]
  _GGMUX2 #(8, 8) g4 (.I0(w121), .I1(w5), .S(fdbk60), .Z(w112));   //: @(-588,1108) /sn:0 /R:1 /w:[ 0 11 11 0 ] /ss:0 /do:0
  //: joint g1236 (w116) @(479, 1848) /w:[ 6 48 5 -1 ]
  //: LED g531 (w341) @(740,44) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g448 (w340) @(357,326) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g453 (w28) @(600,68) /sn:0 /R:1 /anc:1 /w:[ 49 ] /type:0
  //: LED g58 (w55) @(675,479) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  D_FF g1629 (.D(w82), .CP(w116), .Q(w86), .NQ(w260));   //: @(552, 2217) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>239 Ro0<9 Ro1<1 ]
  //: joint g520 (w341) @(733, 66) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g1288 (w215) @(451,188) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g1522 (w357) @(683, 27) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g630 (w183) @(757,438) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1017 (w207) @(384, 277) /anc:1 /w:[ 13 14 16 -1 ]
  //: LED g238 (w224) @(480,139) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  //: joint g816 (w0) @(462, 314) /anc:1 /w:[ 33 34 -1 36 ]
  //: LED g585 (w287) @(794,340) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1052 (w111) @(799, 176) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g334 (w25) @(547, 268) /anc:1 /w:[ 22 24 21 -1 ]
  //: LED g241 (w224) @(432,116) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g1168 (w356) @(416, 245) /anc:1 /w:[ 29 30 32 -1 ]
  //: joint g1897 (w360) @(85, 1641) /w:[ 1 2 48 -1 ]
  D_FF g1631 (.D(w93), .CP(w116), .Q(w91), .NQ(w262));   //: @(813, 2221) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>231 Ro0<0 Ro1<1 ]
  //: joint g1502 (w357) @(679, 39) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g1521 (w151) @(660,-5) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: joint g265 (w29) @(500, 189) /anc:1 /w:[ 10 -1 9 24 ]
  //: LED g272 (w317) @(512,376) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g476 (w300) @(589, 468) /anc:1 /w:[ 4 6 -1 3 ]
  D_FF g1761 (.D(w332), .CP(w34), .Q(w160), .NQ(w324));   //: @(163, 1047) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>73 Ro0<49 Ro1<1 ]
  //: joint g2030 (w215) @(365, 1216) /w:[ 4 6 -1 3 ]
  //: LED g845 (w120) @(439,21) /sn:0 /R:1 /anc:1 /w:[ 23 ] /type:0
  //: LED g1404 (w71) @(542,347) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: LED g53 (w51) @(826,401) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: joint g747 (w204) @(437, 299) /anc:1 /w:[ 29 30 -1 32 ]
  //: joint g554 (w201) @(500, 325) /anc:1 /w:[ 43 -1 44 46 ]
  //: LED g413 (w27) @(513,248) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g957 (w64) @(579,-33) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g1252 (w171) @(748,218) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1680 (w51) @(1194, 1801) /w:[ 2 4 1 -1 ]
  //: joint g548 (w201) @(453, 396) /anc:1 /w:[ 19 -1 20 22 ]
  //: joint g200 (w274) @(349, 192) /anc:1 /w:[ 9 10 12 -1 ]
  //: LED g1382 (w196) @(568,367) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g1648 (w81) @(1258, 2096) /w:[ -1 2 1 8 ]
  //: LED g546 (w201) @(498,348) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: LED g503 (w87) @(727,22) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g2048 (w35) @(325, 1036) /w:[ 4 6 -1 3 ]
  //: LED g526 (w341) @(731,55) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g799 (w24) @(993, 1655) /w:[ 1 2 8 -1 ]
  //: joint g424 (w32) @(570, 116) /anc:1 /w:[ 14 13 28 -1 ]
  //: LED g1578 (w174) @(809,264) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1936 (w51) @(1292, 984) /w:[ -1 6 8 5 ]
  //: LED g624 (w183) @(726,392) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g457 (w28) @(600,-20) /sn:0 /R:1 /anc:1 /w:[ 23 ] /type:0
  //: joint g881 (w75) @(810, 2089) /w:[ 2 4 1 -1 ]
  D_FF g1893 (.D(w274), .CP(w34), .Q(w215), .NQ(w386));   //: @(162, 1484) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>175 Ro0<49 Ro1<1 ]
  //: joint g1906 (w29) @(108, 598) /w:[ -1 4 30 3 ]
  //: LED g193 (w169) @(776,204) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: LED g1019 (w207) @(358,298) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: LED g1601 (w173) @(824,247) /sn:0 /anc:1 /w:[ 21 ] /type:0
  D_FF g1737 (.D(w228), .CP(w34), .Q(w120), .NQ(w291));   //: @(-165, 1624) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>231 Ro0<13 Ro1<1 ]
  //: joint g1178 (w356) @(341, 266) /anc:1 /w:[ 8 -1 7 46 ]
  //: LED g1402 (w304) @(539,415) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  D_FF g1637 (.D(w100), .CP(w116), .Q(w96), .NQ(w267));   //: @(1139, 2226) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>221 Ro0<9 Ro1<1 ]
  //: joint g939 (w211) @(413, 210) /anc:1 /w:[ 29 30 32 -1 ]
  //: joint g1050 (w111) @(748, 185) /anc:1 /w:[ 39 40 -1 42 ]
  //: LED g1173 (w356) @(379,266) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g82 (w86) @(334,96) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: LED g1975 (w101) @(343,5) /sn:0 /w:[ 0 ] /type:3
  D_FF g1795 (.D(w339), .CP(w34), .Q(w332), .NQ(w351));   //: @(99, 1046) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>75 Ro0<49 Ro1<1 ]
  //: LED g650 (w181) @(705,300) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: SWITCH g1894 (w115) @(301,-73) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:0
  //: joint g1924 (w31) @(1264, 864) /w:[ -1 4 6 3 ]
  //: LED g780 (w339) @(772,51) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: joint g1212 (w174) @(796, 273) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g756 (w296) @(491, 16) /anc:1 /w:[ 23 24 -1 26 ]
  //: LED g1105 (w283) @(465,228) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: LED g738 (w204) @(425,320) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: LED g669 (w202) @(461,362) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g1572 (w177) @(765,271) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: LED g89 (w95) @(472,-54) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  _GGMUX2 #(8, 8) g2 (.I0(w7), .I1(w114), .S(fdbk60), .Z(w18));   //: @(281,1780) /sn:0 /R:2 /w:[ 5 1 15 1 ] /ss:0 /do:0
  //: LED g760 (w296) @(475,16) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  D_FF g1628 (.D(w84), .CP(w116), .Q(w93), .NQ(w257));   //: @(749, 2220) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>233 Ro0<0 Ro1<1 ]
  //: LED g786 (w339) @(814,13) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g388 (w166) @(688, 174) /anc:1 /w:[ 13 14 -1 16 ]
  //: LED g1561 (w173) @(773,238) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g883 (w116) @(541, 1848) /w:[ 8 46 7 -1 ]
  //: joint g2052 (w183) @(317, 996) /w:[ 4 6 -1 3 ]
  //: LED g491 (w300) @(599,405) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g1246 (w171) @(773,221) /sn:0 /anc:1 /w:[ 37 ] /type:0
  D_FF g1750 (.D(w186), .CP(w34), .Q(w314), .NQ(w309));   //: @(-362, 1329) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>139 Ro0<49 Ro1<1 ]
  //: LED g868 (w103) @(755,144) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g288 (w286) @(830, 339) /anc:1 /w:[ 11 -1 12 14 ]
  //: joint g411 (w340) @(381, 299) /anc:1 /w:[ 13 14 -1 16 ]
  //: joint g1403 (w71) @(516, 383) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g887 (w16) @(-578, 848) /w:[ 8 38 7 -1 ]
  //: joint g1520 (w357) @(669, 63) /anc:1 /w:[ 43 44 46 -1 ]
  //: LED g599 (w265) @(431,84) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g102 (w153) @(699, 47) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g1097 (w283) @(427,235) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g873 (w70) @(672, 2087) /w:[ 2 4 1 -1 ]
  //: joint g1803 (w300) @(-47, 1347) /w:[ 46 45 48 -1 ]
  //: LED g381 (w166) @(652,177) /sn:0 /anc:1 /w:[ 27 ] /type:0
  //: LED g1261 (w297) @(582,379) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  D_FF g1738 (.D(w286), .CP(w34), .Q(w287), .NQ(w292));   //: @(99, 1189) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>7 Ro0<49 Ro1<1 ]
  //: LED g824 (w0) @(473,316) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: joint g495 (w116) @(446, 1870) /w:[ -1 2 1 96 ]
  //: LED g180 (w21) @(710,263) /sn:0 /anc:1 /w:[ 0 ] /type:0
  //: LED g1593 (w174) @(746,246) /sn:0 /anc:1 /w:[ 41 ] /type:0
  PosBin60 g2077 (.pos(w252), .bin(w38));   //: @(-93, 477) /sz:(95, 40) /sn:0 /p:[ Li0>1 Ro0<1 ]
  //: LED g547 (w201) @(482,372) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g1499 (w357) @(673, 51) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g168 (w21) @(662,239) /sn:0 /anc:1 /w:[ 27 ] /type:0
  //: LED g1412 (w71) @(499,457) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: LED g1316 (w134) @(616,43) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: LED g1128 (w108) @(565,18) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g565 (w201) @(521,316) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g1474 (w219) @(364,133) /sn:0 /R:2 /anc:1 /w:[ 17 ] /type:0
  //: comment g1990 @(298,186)
  //: /line:"<h1 color=blue>9</h1>"
  //: /end
  //: joint g518 (w87) @(762, -14) /anc:1 /w:[ 7 -1 8 10 ]
  //: joint g2024 (w228) @(382, 1276) /w:[ 6 8 -1 5 ]
  //: joint g282 (w317) @(511, 340) /anc:1 /w:[ 43 -1 44 46 ]
  assign w252 = {w64, w108, w141, w360, w233, w296, w120, w228, w265, w224, w290, w219, w352, w215, w274, w211, w283, w356, w207, w340, w204, w0, w202, w201, w317, w71, w304, w196, w297, w300, w33, w35, w113, w314, w186, w183, w298, w181, w287, w286, w177, w174, w173, w171, w169, w89, w111, w330, w103, w160, w332, w339, w341, w87, w153, w357, w151, w163, w134, w28}; //: CONCAT g2016  @(552,1051) /sn:0 /w:[ 0 5 0 0 5 7 7 7 7 5 5 5 7 7 5 5 5 5 5 0 5 5 5 5 5 5 5 0 5 5 0 5 5 0 5 5 5 5 5 5 5 5 0 5 5 5 0 0 5 0 5 5 5 5 0 5 5 5 5 5 7 ] /dr:1 /tp:0 /drp:1
  //: LED g754 (w296) @(506,63) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: LED g559 (w201) @(459,408) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1463 (w290) @(422, 119) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1208 (w151) @(646,45) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1804 (w332) @(148, 1060) /w:[ 1 2 48 -1 ]
  //: joint g974 (w103) @(755, 154) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g1425 (w196) @(556,430) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g1921 (w14) @(1256, 824) /w:[ -1 2 1 4 ]
  //: LED g684 (w228) @(463,81) /sn:0 /R:2 /anc:1 /w:[ 37 ] /type:0
  //: joint g1306 (w134) @(633, -20) /anc:1 /w:[ -1 19 20 22 ]
  //: LED g644 (w181) @(737,327) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g366 (w233) @(516, 8) /anc:1 /w:[ 23 24 -1 26 ]
  //: joint g1028 (w207) @(371, 283) /anc:1 /w:[ 9 10 12 -1 ]
  //: joint g1656 (w73) @(929, 1797) /w:[ 6 5 8 -1 ]
  //: frame g1995 @(256,-114) /sn:0 /wi:649 /ht:624 /tx:"Analog  clock"
  //: joint g1933 (w47) @(1286, 954) /w:[ -1 6 8 5 ]
  //: joint g1947 (w62) @(1318, 1094) /w:[ -1 4 6 3 ]
  //: LED g666 (w202) @(452,373) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g955 (w64) @(580,-20) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g913 (w33) @(613,354) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g450 (w340) @(369, 304) /anc:1 /w:[ 9 10 -1 12 ]
  //: joint g1349 (w116) @(540, 1995) /w:[ 102 140 101 -1 ]
  //: LED g254 (w29) @(525,202) /sn:0 /R:2 /anc:1 /w:[ 21 ] /type:0
  //: LED g860 (w207) @(445,262) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g1134 (w330) @(847, 142) /anc:1 /w:[ 11 12 14 -1 ]
  D_FF g1335 (.D(w48), .CP(w116), .Q(w50), .NQ(w178));   //: @(1077, 1786) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>31 Ro0<0 Ro1<1 ]
  //: joint g620 (w183) @(710, 392) /anc:1 /w:[ 23 24 -1 26 ]
  //: LED g1501 (w163) @(631,43) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1175 (w356) @(379, 256) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g891 (w33) @(607, 404) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1061 (w111) @(773, 181) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1818 (w317) @(280, 1352) /w:[ -1 2 1 48 ]
  //: joint g419 (w32) @(582, 140) /anc:1 /w:[ 20 19 26 -1 ]
  //: joint g1384 (w196) @(551, 391) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g115 (w20) @(600,81) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g1428 (w71) @(507, 408) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1301 (w215) @(349, 166) /anc:1 /w:[ 9 10 12 -1 ]
  //: LED g75 (w76) @(327,281) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: joint g1269 (w297) @(569, 391) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g777 (w339) @(804, 35) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g39 (w9) @(739, 1651) /w:[ 2 4 1 -1 ]
  //: LED g1532 (w151) @(672,-44) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g1110 (w108) @(582, 56) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1081 (w35) @(621, 378) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1721 (w174) @(-49, 1200) /w:[ 46 45 48 -1 ]
  //: joint g673 (w228) @(397, 16) /anc:1 /w:[ 11 -1 12 14 ]
  //: joint g1016 (w207) @(358, 288) /anc:1 /w:[ 5 6 8 -1 ]
  //: LED g485 (w300) @(599,468) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g455 (w28) @(610, -58) /anc:1 /w:[ -1 9 10 12 ]
  //: LED g1176 (w356) @(429,251) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: LED g1300 (w215) @(362,179) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1570 (w174) @(783, 270) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1701 (w34) @(-113, 1690) /w:[ 210 228 209 -1 ]
  //: LED g201 (w169) @(864,204) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g700 (w332) @(811, 76) /anc:1 /w:[ 15 16 -1 18 ]
  //: LED g1487 (w352) @(464,176) /sn:0 /R:2 /anc:1 /w:[ 49 ] /type:0
  //: joint g1638 (w116) @(477, 2287) /w:[ 198 240 197 -1 ]
  //: joint g1880 (w89) @(-307, 1196) /w:[ 46 45 48 -1 ]
  //: joint g966 (w64) @(594, 30) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1681 (w63) @(1197, 1948) /w:[ 1 2 8 -1 ]
  D_FF g1227 (.D(w27), .CP(w16), .Q(w29), .NQ(w139));   //: @(-174, 786) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>27 Ro0<33 Ro1<1 ]
  //: joint g236 (w224) @(372, 69) /anc:1 /w:[ 10 9 -1 44 ]
  //: LED g908 (w89) @(764,189) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: LED g488 (w300) @(599,417) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g1635 (w116) @(930, 2287) /w:[ 212 226 211 -1 ]
  //: LED g832 (w120) @(497,86) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g316 (w25) @(555, 256) /anc:1 /w:[ 26 28 25 -1 ]
  //: joint g1910 (w22) @(100, 638) /w:[ -1 25 26 28 ]
  //: comment g1984 @(887,193)
  //: /line:"<h1 color=blue>3</h1>"
  //: /end
  //: joint g1861 (w0) @(-306, 1490) /w:[ 1 2 48 -1 ]
  D_FF g1745 (.D(w181), .CP(w34), .Q(w298), .NQ(w299));   //: @(226, 1191) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 Ro1<1 ]
  //: joint g1163 (w113) @(648, 413) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g1806 (w34) @(-239, 1545) /w:[ 156 186 155 -1 ]
  //: LED g688 (w228) @(474,90) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  //: joint g2049 (w113) @(323, 1026) /w:[ 1 2 -1 44 ]
  //: joint g558 (w201) @(439, 420) /anc:1 /w:[ 11 -1 12 14 ]
  //: frame g1997 @(-777,712) /sn:0 /wi:799 /ht:160 /tx:"sequence of flip-flops as shift register"
  //: joint g3 (fdbk60) @(236, 1755) /w:[ 14 -1 13 16 ]
  //: LED g1071 (w35) @(644,442) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1960 (w77) @(1347, 1224) /w:[ -1 6 8 5 ]
  //: LED g542 (w181) @(814,390) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: LED g373 (w340) @(417,296) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g1124 (w108) @(571, -7) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g962 (w64) @(590, -20) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g1255 (w171) @(824,225) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1902 (w166) @(94, 668) /w:[ -1 4 30 3 ]
  //: joint g183 (w169) @(788, 216) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1025 (w207) @(396, 272) /anc:1 /w:[ 17 18 20 -1 ]
  D_FF g1345 (.D(w54), .CP(w116), .Q(w53), .NQ(w210));   //: @(553, 1925) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>141 Ro0<9 Ro1<1 ]
  //: joint g940 (w211) @(362, 214) /anc:1 /w:[ 13 14 16 -1 ]
  //: LED g129 (w153) @(717,-25) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g1364 (w52) @(1259, 1802) /w:[ -1 2 8 1 ]
  //: joint g2066 (w160) @(279, 856) /w:[ 4 6 -1 3 ]
  //: joint g1811 (w34) @(-112, 1545) /w:[ 160 182 159 -1 ]
  //: LED g305 (w286) @(782,298) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g1239 (w171) @(862,230) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g1550 (w174) @(746, 258) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1886 (w34) @(-438, 1545) /w:[ 150 192 149 -1 ]
  D_FF g1889 (.D(w352), .CP(w34), .Q(w219), .NQ(w384));   //: @(-490, 1619) /sz:(40, 56) /sn:0 /p:[ Li0>13 Li1>241 Ro0<0 Ro1<1 ]
  //: joint g1274 (w297) @(570, 379) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g1386 (w196) @(559,417) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1775 (w171) @(-175, 1198) /w:[ 1 2 48 -1 ]
  //: joint g580 (w287) @(758, 330) /anc:1 /w:[ 31 -1 32 34 ]
  //: LED g811 (w0) @(388,393) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g705 (w332) @(811,63) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g680 (w228) @(386, 7) /anc:1 /w:[ 10 9 -1 48 ]
  //: LED g459 (w28) @(600,18) /sn:0 /R:1 /anc:1 /w:[ 35 ] /type:0
  //: LED g67 (w65) @(470,462) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g602 (w265) @(431, 71) /anc:1 /w:[ 25 -1 26 28 ]
  //: joint g2059 (w173) @(299, 926) /w:[ 4 6 -1 3 ]
  //: joint g1837 (w34) @(88, 1251) /w:[ 5 6 8 -1 ]
  //: LED g257 (w224) @(444,121) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: joint g1651 (w42) @(608, 1792) /w:[ 6 5 8 -1 ]
  //: joint g1938 (w54) @(1300, 1004) /w:[ -1 4 6 3 ]
  //: LED g350 (w67) @(516,157) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g109 (w19) @(713,204) /sn:0 /anc:1 /w:[ 9 ] /type:0
  _GGOR2 #(6) g1719 (.I0(w104), .I1(w26), .Z(w16));   //: @(-801,641) /sn:0 /w:[ 0 1 0 ]
  //: LED g264 (w29) @(487,202) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: LED g56 (w53) @(729,461) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g805 (w116) @(867, 1705) /w:[ 64 82 63 -1 ]
  //: joint g1780 (w340) @(-168, 1492) /w:[ 1 2 48 -1 ]
  //: joint g735 (w204) @(449, 293) /anc:1 /w:[ 33 34 -1 36 ]
  //: joint g1055 (w111) @(850, 166) /anc:1 /w:[ 7 8 10 -1 ]
  D_FF g1768 (.D(w108), .CP(w34), .Q(w64), .NQ(w336));   //: @(224, 1630) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>219 Ro0<0 Ro1<1 ]
  //: joint g733 (w204) @(402, 321) /anc:1 /w:[ 17 18 -1 20 ]
  //: joint g682 (w228) @(408, 24) /anc:1 /w:[ 15 -1 16 18 ]
  //: joint g1560 (w173) @(785, 252) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g333 (w25) @(559,280) /sn:0 /R:3 /anc:1 /w:[ 19 ] /type:0
  //: joint g1352 (w116) @(605, 1995) /w:[ 104 138 103 -1 ]
  //: joint g1608 (w116) @(540, 2142) /w:[ 150 192 149 -1 ]
  //: joint g2026 (w224) @(378, 1256) /w:[ 4 6 -1 3 ]
  //: joint g1650 (w132) @(543, 1791) /w:[ 1 2 8 -1 ]
  //: LED g649 (w181) @(759,345) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g1151 (w113) @(645, 401) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g583 (w287) @(734, 313) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g283 (w317) @(506, 352) /anc:1 /w:[ 39 -1 40 42 ]
  //: LED g1289 (w215) @(388,182) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g242 (w224) @(444, 104) /anc:1 /w:[ 29 -1 30 32 ]
  //: LED g281 (w317) @(517,364) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g1943 (w57) @(1310, 1054) /w:[ -1 4 6 3 ]
  //: joint g1711 (w22) @(-385, 796) /w:[ 30 29 32 -1 ]
  //: LED g675 (w228) @(397,27) /sn:0 /R:2 /anc:1 /w:[ 13 ] /type:0
  //: joint g422 (w32) @(587, 152) /anc:1 /w:[ 22 21 24 -1 ]
  //: LED g1379 (w71) @(503,445) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g157 (w21) @(686, 269) /anc:1 /w:[ -1 18 20 17 ]
  //: LED g324 (w186) @(680,363) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g1939 (w53) @(1302, 1014) /w:[ -1 4 6 3 ]
  //: LED g721 (w298) @(742,367) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g785 (w339) @(794, 44) /anc:1 /w:[ 15 16 -1 18 ]
  //: joint g1045 (w360) @(531, 0) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1460 (w352) @(349,154) /sn:0 /R:2 /anc:1 /w:[ 0 ] /type:0
  //: LED g617 (w265) @(487,123) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g166 (w21) @(698,257) /sn:0 /anc:1 /w:[ 15 ] /type:0
  //: LED g1319 (w134) @(618,19) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: LED g365 (w233) @(489,-16) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g1415 (w196) @(561,404) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g28 (w19) @(663, 221) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g522 (w183) @(680,321) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g536 (w341) @(758,22) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g464 (w28) @(600,-58) /sn:0 /R:1 /anc:1 /w:[ 11 ] /type:0
  //: joint g938 (w211) @(437, 208) /anc:1 /w:[ 37 38 40 -1 ]
  //: joint g1539 (w151) @(686, -56) /anc:1 /w:[ -1 7 8 10 ]
  //: joint g1323 (w134) @(632, -7) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1511 (w357) @(676,15) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  D_FF g1649 (.D(w91), .CP(w116), .Q(w90), .NQ(w276));   //: @(876, 2222) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>229 Ro0<0 Ro1<1 ]
  D_FF g888 (.D(w29), .CP(w16), .Q(w67), .NQ(w125));   //: @(-110, 787) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>25 Ro0<33 Ro1<1 ]
  //: joint g1000 (w314) @(688, 458) /anc:1 /w:[ 8 10 -1 7 ]
  //: joint g296 (w286) @(794, 322) /anc:1 /w:[ 23 -1 24 26 ]
  //: LED g1543 (w151) @(664,-18) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g1555 (w177) @(839,300) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g1923 (w12) @(1260, 844) /w:[ -1 4 6 3 ]
  //: joint g925 (w33) @(611, 455) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g1495 (w151) @(639,71) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: LED g964 (w64) @(583,18) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g1251 (w171) @(773, 233) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g601 (w265) @(455, 87) /anc:1 /w:[ 33 -1 34 36 ]
  //: LED g1375 (w71) @(538,359) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g1577 (w177) @(741, 273) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1914 (w5) @(1244, 764) /w:[ -1 6 8 5 ]
  //: joint g515 (w87) @(708, 70) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g1260 (w297) @(578,430) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g80 (w81) @(323,147) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: joint g1677 (w80) @(1062, 2093) /w:[ 1 2 8 -1 ]
  D_FF g1778 (.D(w341), .CP(w34), .Q(w339), .NQ(w342));   //: @(33, 1045) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>77 Ro0<49 Ro1<1 ]
  D_FF g1868 (.D(w224), .CP(w34), .Q(w265), .NQ(w381));   //: @(-295, 1622) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>235 Ro0<49 Ro1<1 ]
  D_FF g1757 (.D(w314), .CP(w34), .Q(w113), .NQ(w320));   //: @(-294, 1330) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>137 Ro0<49 Ro1<1 ]
  D_FF g810 (.D(w12), .CP(w116), .Q(w11), .NQ(w49));   //: @(1077, 1643) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>77 Ro0<0 Ro1<1 ]
  //: LED g291 (w286) @(794,304) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g510 (w87) @(735,10) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g379 (w340) @(453, 263) /anc:1 /w:[ 37 38 -1 40 ]
  //: joint g1468 (w219) @(440, 144) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1905 (w25) @(104, 618) /w:[ -1 4 30 3 ]
  //: joint g693 (w332) @(833, 60) /anc:1 /w:[ 7 8 -1 10 ]
  //: LED g613 (w265) @(371,46) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g198 (w169) @(852, 216) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g51 (w19) @(663,204) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: joint g662 (w202) @(422, 395) /anc:1 /w:[ 15 -1 16 18 ]
  //: joint g519 (w87) @(769, -26) /anc:1 /w:[ -1 3 4 6 ]
  //: LED g302 (w286) @(758,287) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g804 (w14) @(928, 1654) /w:[ 6 5 8 -1 ]
  //: joint g538 (w341) @(779, 11) /anc:1 /w:[ 15 -1 16 18 ]
  //: LED g290 (w286) @(722,269) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: LED g460 (w28) @(600,-46) /sn:0 /R:1 /anc:1 /w:[ 15 ] /type:0
  //: joint g1418 (w304) @(527, 415) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g72 (w75) @(344,334) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: LED g182 (w21) @(686,251) /sn:0 /anc:1 /w:[ 19 ] /type:0
  //: joint g1782 (w34) @(-501, 1690) /w:[ 198 240 197 -1 ]
  //: LED g1139 (w330) @(746,162) /sn:0 /anc:1 /w:[ 45 ] /type:0
  D_FF g1365 (.D(w57), .CP(w116), .Q(w58), .NQ(w226));   //: @(877, 1930) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>131 Ro0<9 Ro1<1 ]
  //: joint g545 (w201) @(460, 384) /anc:1 /w:[ 23 -1 24 26 ]
  //: joint g657 (w202) @(440, 373) /anc:1 /w:[ 23 -1 24 26 ]
  //: joint g444 (w340) @(405, 287) /anc:1 /w:[ 21 22 -1 24 ]
  //: LED g840 (w120) @(459,42) /sn:0 /R:1 /anc:1 /w:[ 31 ] /type:0
  //: LED g570 (w332) @(776,86) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g2065 (w103) @(281, 866) /w:[ 1 2 -1 44 ]
  //: LED g187 (w169) @(826,204) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1716 (w41) @(-321, 797) /w:[ 1 2 32 -1 ]
  //: joint g619 (w183) @(691, 357) /anc:1 /w:[ 35 36 -1 38 ]
  //: LED g348 (w67) @(552,175) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: LED g1083 (w35) @(638,416) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1840 (w283) @(17, 1495) /w:[ 1 2 48 -1 ]
  //: LED g1472 (w290) @(348,102) /sn:0 /R:2 /anc:1 /w:[ 9 ] /type:0
  //: joint g914 (w33) @(608, 416) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1166 (w113) @(656, 439) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g751 (w204) @(368, 346) /anc:1 /w:[ -1 8 7 46 ]
  //: joint g2025 (w265) @(380, 1266) /w:[ 4 6 -1 3 ]
  //: joint g894 (w89) @(813, 195) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g1121 (w108) @(578, 31) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g145 (w160) @(736,135) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1226 (w16) @(-645, 848) /w:[ 6 40 5 -1 ]
  //: joint g608 (w265) @(371, 34) /anc:1 /w:[ 8 7 -1 46 ]
  //: joint g407 (w27) @(537, 221) /anc:1 /w:[ -1 18 17 24 ]
  //: LED g1406 (w196) @(553,443) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: LED g911 (w33) @(622,467) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1784 (w224) @(-308, 1635) /w:[ 1 2 48 -1 ]
  //: joint g2067 (w332) @(277, 846) /w:[ 4 6 -1 3 ]
  //: joint g1042 (w360) @(546, 37) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1858 (w34) @(215, 1545) /w:[ 170 172 169 -1 ]
  //: joint g1652 (w156) @(671, 1793) /w:[ 6 5 8 -1 ]
  D_FF g1766 (.D(w169), .CP(w34), .Q(w171), .NQ(w331));   //: @(-227, 1184) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>27 Ro0<49 Ro1<1 ]
  //: joint g351 (w67) @(516, 139) /anc:1 /w:[ -1 10 12 9 ]
  //: LED g125 (w153) @(705,-1) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  D_FF g1221 (.D(w25), .CP(w16), .Q(w27), .NQ(w129));   //: @(-240, 785) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>29 Ro0<33 Ro1<1 ]
  D_FF g806 (.D(w3), .CP(w116), .Q(w6), .NQ(w99));   //: @(617, 1636) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>91 Ro0<9 Ro1<1 ]
  //: joint g632 (w183) @(684, 345) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1907 (w32) @(112, 578) /w:[ -1 6 32 5 ]
  //: joint g275 (w317) @(482, 400) /anc:1 /w:[ 23 -1 24 26 ]
  D_FF g1353 (.D(w62), .CP(w116), .Q(w63), .NQ(w217));   //: @(1140, 1934) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>123 Ro0<9 Ro1<1 ]
  //: joint g1770 (w34) @(19, 1690) /w:[ 214 224 213 -1 ]
  //: LED g1517 (w151) @(651,33) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g1955 (w74) @(1337, 1174) /w:[ -1 4 6 3 ]
  //: joint g279 (w317) @(470, 424) /anc:1 /w:[ 15 -1 16 18 ]
  //: joint g579 (w287) @(806, 360) /anc:1 /w:[ 15 -1 16 18 ]
  //: joint g1431 (w219) @(403, 133) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1264 (w297) @(585,354) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g783 (w339) @(718, 110) /anc:1 /w:[ 43 44 -1 46 ]
  //: joint g1952 (w70) @(1331, 1144) /w:[ -1 6 8 5 ]
  //: LED g719 (w298) @(695,312) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g352 (w67) @(564,181) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g1496 (w163) @(628,56) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g725 (w298) @(714,334) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g1588 (w177) @(851,304) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: LED g1009 (w314) @(668,384) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g1525 (w163) @(646,-33) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  D_FF g1792 (.D(w211), .CP(w34), .Q(w274), .NQ(w349));   //: @(98, 1483) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>177 Ro0<49 Ro1<1 ]
  //: joint g1965 (w84) @(1360, 1274) /w:[ -1 4 6 3 ]
  //: LED g1452 (w290) @(410,126) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: LED g1077 (w35) @(631,378) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g1678 (w48) @(1067, 1799) /w:[ 2 4 1 -1 ]
  //: joint g1765 (w215) @(213, 1498) /w:[ 1 2 48 -1 ]
  //: joint g997 (w314) @(673, 421) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g442 (w340) @(441,284) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g555 (w201) @(493, 336) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g150 (w160) @(748, 144) /anc:1 /w:[ 39 40 -1 42 ]
  //: LED g1453 (w290) @(397,122) /sn:0 /R:2 /anc:1 /w:[ 21 ] /type:0
  //: LED g481 (w300) @(599,456) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g447 (w340) @(393, 294) /anc:1 /w:[ 17 18 -1 20 ]
  //: joint g714 (w298) @(749, 388) /anc:1 /w:[ 19 20 -1 22 ]
  //: LED g897 (w89) @(839,183) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g1278 (w297) @(580,404) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g1051 (w111) @(837,158) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g833 (w120) @(452, 21) /anc:1 /w:[ 21 22 -1 24 ]
  D_FF g1348 (.D(w56), .CP(w116), .Q(w55), .NQ(w214));   //: @(684, 1927) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>137 Ro0<9 Ro1<1 ]
  //: joint g1755 (w181) @(216, 1204) /w:[ 1 2 48 -1 ]
  //: joint g1604 (w177) @(802, 296) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1466 (w352) @(362,156) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: joint g1186 (w356) @(366, 260) /anc:1 /w:[ 13 14 16 -1 ]
  //: joint g1374 (w304) @(545, 352) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g1326 (w134) @(619,6) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g948 (w211) @(437,218) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  D_FF g875 (.D(w156), .CP(w116), .Q(w40), .NQ(w172));   //: @(685, 1780) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>43 Ro0<0 Ro1<1 ]
  //: joint g1726 (w34) @(-177, 1545) /w:[ 158 184 157 -1 ]
  //: joint g1076 (w35) @(631, 429) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g722 (w298) @(778, 419) /anc:1 /w:[ 8 -1 10 7 ]
  //: joint g1665 (w54) @(543, 1938) /w:[ 1 2 8 -1 ]
  D_FF g1756 (.D(w207), .CP(w34), .Q(w356), .NQ(w318));   //: @(-101, 1480) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>183 Ro0<49 Ro1<1 ]
  //: LED g1215 (w171) @(785,222) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g483 (w300) @(589, 368) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1277 (w297) @(563, 456) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g473 (w300) @(599,443) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g1102 (w283) @(338,252) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g549 (w201) @(485, 348) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g44 (w46) @(876,257) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g935 (w211) @(375,223) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: joint g681 (w228) @(485, 87) /anc:1 /w:[ 43 -1 44 46 ]
  _GGMUX2 #(8, 8) g1663 (.I0(w8), .I1(w32), .S(fdbk60), .Z(w109));   //: @(-868,791) /sn:0 /R:1 /w:[ 1 3 7 1 ] /ss:0 /do:0
  //: LED g54 (w52) @(801,431) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: LED g40 (w40) @(878,204) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g1015 (w207) @(384,287) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1819 (w34) @(-47, 1545) /w:[ 162 180 161 -1 ]
  D_FF g1824 (.D(w265), .CP(w34), .Q(w228), .NQ(w365));   //: @(-229, 1623) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>233 Ro0<0 Ro1<1 ]
  //: LED g1424 (w304) @(535,428) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1708 (w166) @(-582, 793) /w:[ 1 2 32 -1 ]
  //: joint g2055 (w287) @(307, 966) /w:[ 4 6 -1 3 ]
  //: joint g1617 (w116) @(866, 2142) /w:[ 160 182 159 -1 ]
  //: joint g1587 (w173) @(748, 244) /anc:1 /w:[ 43 44 46 -1 ]
  //: LED g1562 (w173) @(811,244) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: joint g506 (w87) @(716, 58) /anc:1 /w:[ 31 -1 32 34 ]
  //: joint g1895 (w103) @(281, 1062) /w:[ -1 45 46 48 ]
  //: joint g1563 (w173) @(773, 250) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g462 (w28) @(610, 42) /anc:1 /w:[ 41 42 44 -1 ]
  //: joint g1670 (w57) @(866, 1943) /w:[ 1 2 8 -1 ]
  //: LED g65 (w62) @(518,480) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: frame g1998 @(440,1616) /sn:0 /wi:860 /ht:700 /tx:"sequence of flip-flops as shift register"
  //: LED g1144 (w330) @(733,166) /sn:0 /anc:1 /w:[ 47 ] /type:0
  D_FF g1234 (.D(w132), .CP(w116), .Q(w42), .NQ(w168));   //: @(554, 1778) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>47 Ro0<9 Ro1<1 ]
  //: joint g304 (w286) @(746, 298) /anc:1 /w:[ -1 40 42 39 ]
  //: joint g634 (w183) @(704, 381) /anc:1 /w:[ 27 28 -1 30 ]
  //: LED g1078 (w35) @(646,455) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g1342 (w116) @(1065, 1995) /w:[ 118 124 117 -1 ]
  //: joint g2041 (w317) @(339, 1106) /w:[ 4 6 -1 3 ]
  //: LED g863 (w141) @(555,45) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g427 (w32) @(565, 104) /anc:1 /w:[ 12 11 30 -1 ]
  //: LED g686 (w228) @(430,54) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: joint g1609 (w116) @(998, 2142) /w:[ 164 178 163 -1 ]
  //: joint g1833 (w228) @(-176, 1637) /w:[ 2 4 1 -1 ]
  //: comment g1982 @(280,-63) /sn:0
  //: /line:"<h3 color=blue>+1 m</h3>"
  //: /end
  //: joint g1860 (w27) @(-187, 799) /w:[ 1 2 32 -1 ]
  //: joint g245 (w224) @(408, 86) /anc:1 /w:[ 17 -1 18 20 ]
  //: joint g1090 (w283) @(452, 221) /anc:1 /w:[ 41 42 -1 44 ]
  //: LED g564 (w201) @(451,420) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g1202 (w141) @(541,-4) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g1643 (w116) @(738, 2287) /w:[ 206 232 205 -1 ]
  //: LED g1417 (w304) @(557,352) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g131 (w20) @(600,156) /sn:0 /R:1 /anc:1 /w:[ 31 ] /type:0
  //: LED g1004 (w314) @(678,409) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g690 (w228) @(495,108) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g1481 (w290) @(422,131) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: joint g1229 (w116) @(606, 1848) /w:[ 10 44 9 -1 ]
  //: LED g727 (w298) @(723,345) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: LED g1167 (w113) @(651,389) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g598 (w265) @(455,100) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g1224 (w16) @(-384, 848) /w:[ 14 32 13 -1 ]
  //: LED g1321 (w134) @(613,69) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: LED g1043 (w360) @(500,-49) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g1862 (w29) @(-122, 800) /w:[ 1 2 32 -1 ]
  //: joint g1626 (w116) @(1064, 2287) /w:[ 216 222 215 -1 ]
  D_FF g874 (.D(w67), .CP(w16), .Q(w32), .NQ(w118));   //: @(-47, 788) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>23 Ro0<0 Ro1<1 ]
  //: joint g347 (w233) @(495, -40) /anc:1 /w:[ 10 9 48 -1 ]
  //: joint g890 (w103) @(779, 144) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1315 (w134) @(638, -58) /anc:1 /w:[ -1 7 8 10 ]
  //: LED g60 (w32) @(543,92) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: LED g210 (w41) @(599,254) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g1928 (w156) @(1276, 904) /w:[ -1 2 1 4 ]
  //: joint g2072 (w357) @(267, 796) /w:[ 4 6 -1 3 ]
  //: joint g1422 (w196) @(537, 468) /anc:1 /w:[ 8 10 -1 7 ]
  //: joint g126 (w153) @(723, -1) /anc:1 /w:[ 19 -1 20 22 ]
  //: joint g185 (w169) @(751, 216) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1724 (w286) @(89, 1202) /w:[ 1 2 48 -1 ]
  //: joint g1483 (w290) @(385, 105) /anc:1 /w:[ 18 -1 17 44 ]
  //: LED g593 (w287) @(714,285) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: joint g1457 (w352) @(375, 147) /anc:1 /w:[ 21 22 24 -1 ]
  //: joint g1258 (w297) @(566, 430) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g946 (w211) @(425, 209) /anc:1 /w:[ 33 34 36 -1 ]
  //: joint g1735 (w34) @(-46, 1251) /w:[ 13 14 16 -1 ]
  //: joint g1865 (w34) @(-532, 1545) /w:[ 146 145 -1 196 ]
  //: LED g1250 (w171) @(837,227) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g1969 (w95) @(1368, 1314) /w:[ -1 6 8 5 ]
  //: joint g776 (w339) @(772, 63) /anc:1 /w:[ 23 24 -1 26 ]
  //: joint g691 (w228) @(419, 32) /anc:1 /w:[ 19 -1 20 22 ]
  //: LED g999 (w314) @(694,447) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g1497 (w357) @(701, -23) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g900 (w89) @(839, 193) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g1119 (w108) @(562, -58) /anc:1 /w:[ -1 3 4 6 ]
  //: joint g1109 (w108) @(575, 18) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g112 (w19) @(688, 221) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g689 (w228) @(441,63) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: LED g1582 (w173) @(837,250) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g1193 (w141) @(537,-17) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  D_FF g1823 (.D(w171), .CP(w34), .Q(w173), .NQ(w364));   //: @(-163, 1185) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>23 Ro0<49 Ro1<1 ]
  //: joint g1796 (w25) @(-256, 798) /w:[ 1 2 32 -1 ]
  //: joint g867 (w330) @(784, 161) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g64 (w60) @(544,483) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: LED g263 (w317) @(488,424) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g259 (w224) @(468, 115) /anc:1 /w:[ 37 -1 38 40 ]
  //: joint g540 (w341) @(716, 88) /anc:1 /w:[ 43 -1 44 46 ]
  //: joint g1810 (w34) @(-112, 1398) /w:[ 112 130 111 -1 ]
  //: joint g1867 (w204) @(-243, 1491) /w:[ 1 2 48 -1 ]
  //: LED g676 (w228) @(485,99) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g819 (w0) @(473, 305) /anc:1 /w:[ 37 38 -1 40 ]
  //: LED g1312 (w134) @(614,56) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g609 (w265) @(407,68) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: joint g2020 (w360) @(390, 1316) /w:[ 4 6 -1 3 ]
  //: joint g1900 (w34) @(-238, 1251) /w:[ 25 26 28 -1 ]
  //: LED g1273 (w297) @(586,341) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: joint g1143 (w330) @(808, 154) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g713 (w298) @(704,323) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: LED g843 (w120) @(468,53) /sn:0 /R:1 /anc:1 /w:[ 35 ] /type:0
  //: joint g1657 (w47) @(998, 1798) /w:[ 2 4 1 -1 ]
  //: LED g1473 (w219) @(351,130) /sn:0 /R:2 /anc:1 /w:[ 13 ] /type:0
  //: joint g821 (w0) @(388, 380) /anc:1 /w:[ -1 8 7 46 ]
  D_FF g1347 (.D(w69), .CP(w116), .Q(w57), .NQ(w212));   //: @(814, 1929) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>133 Ro0<9 Ro1<1 ]
  //: LED g1540 (w357) @(671,27) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g1203 (w141) @(551, -4) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g1039 (w360) @(505,-38) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g861 (w211) @(400, 211) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g1093 (w283) @(439, 223) /anc:1 /w:[ 37 38 40 -1 ]
  //: joint g582 (w287) @(723, 306) /anc:1 /w:[ 43 -1 44 46 ]
  //: joint g301 (w286) @(806, 328) /anc:1 /w:[ 19 -1 20 22 ]
  //: LED g207 (w169) @(852,204) /sn:0 /anc:1 /w:[ 13 ] /type:0
  D_FF g1885 (.D(w134), .CP(w34), .Q(w163), .NQ(w383));   //: @(-361, 1039) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>89 Ro0<49 Ro1<1 ]
  //: joint g1378 (w71) @(498, 433) /anc:1 /w:[ 15 16 18 -1 ]
  D_FF g1751 (.D(w204), .CP(w34), .Q(w340), .NQ(w311));   //: @(-228, 1478) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>187 Ro0<49 Ro1<1 ]
  D_FF g1849 (.D(w160), .CP(w34), .Q(w103), .NQ(w377));   //: @(226, 1048) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>71 Ro0<47 Ro1<1 ]
  //: joint g29 (fdbk60) @(-616, 1151) /w:[ 10 9 -1 12 ]
  //: LED g1065 (w111) @(735,178) /sn:0 /anc:1 /w:[ 43 ] /type:0
  //: joint g1967 (w91) @(1364, 1294) /w:[ -1 6 8 5 ]
  //: LED g1213 (w171) @(761,220) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g106 (w153) @(676,59) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1248 (w171) @(761, 232) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g174 (w160) @(820,93) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g494 (w298) @(753,377) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g402 (w22) @(620,243) /sn:0 /R:3 /anc:1 /w:[ 23 ] /type:0
  //: LED g516 (w87) @(719,34) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: joint g1625 (w116) @(800, 2287) /w:[ 208 230 207 -1 ]
  //: joint g1440 (w290) @(446, 129) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g375 (w340) @(357, 308) /anc:1 /w:[ -1 8 7 46 ]
  //: LED g1320 (w134) @(624,-46) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g21 (w14) @(766,-39) /sn:0 /R:1 /anc:1 /w:[ 3 ] /type:0
  //: LED g172 (w160) @(808,99) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g836 (w120) @(489, 64) /anc:1 /w:[ 37 38 -1 40 ]
  //: LED g1088 (w35) @(634,391) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g487 (w300) @(599,380) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g256 (w224) @(396, 80) /anc:1 /w:[ 13 -1 14 16 ]
  //: joint g141 (w153) @(709, 23) /anc:1 /w:[ 27 -1 28 30 ]
  //: LED g341 (w67) @(540,169) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: joint g386 (w166) @(652, 191) /anc:1 /w:[ 25 26 -1 28 ]
  //: LED g222 (w274) @(337,202) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g492 (w300) @(599,368) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g635 (w183) @(744, 438) /anc:1 /w:[ 8 -1 10 7 ]
  //: joint g1671 (w58) @(931, 1944) /w:[ 1 2 8 -1 ]
  //: joint g1908 (w67) @(110, 588) /w:[ -1 4 30 3 ]
  //: LED g562 (w201) @(505,336) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g968 (w64) @(585,42) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1777 (w34) @(-178, 1690) /w:[ 208 230 207 -1 ]
  //: joint g1148 (w113) @(641, 389) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g49 (w48) @(856,334) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g858 (w283) @(439,233) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: LED g137 (w153) @(711,-13) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g1504 (w163) @(634,31) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g953 (w64) @(586,55) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g1285 (w215) @(426,185) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g217 (w274) @(388, 192) /anc:1 /w:[ 21 22 24 -1 ]
  //: joint g1664 (w76) @(929, 2091) /w:[ 1 2 8 -1 ]
  //: joint g2056 (w286) @(305, 956) /w:[ 4 6 -1 3 ]
  //: LED g557 (w201) @(466,396) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g1614 (w116) @(1127, 2142) /w:[ 168 174 167 -1 ]
  //: LED g646 (w181) @(770,354) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: joint g1243 (w171) @(824, 237) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g642 (w181) @(792, 384) /anc:1 /w:[ 15 -1 16 18 ]
  //: LED g628 (w183) @(702,357) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g916 (w33) @(603, 354) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1848 (w160) @(214, 1061) /w:[ 1 2 48 -1 ]
  //: joint g878 (w116) @(932, 1705) /w:[ 66 80 65 -1 ]
  //: LED g420 (w32) @(549,104) /sn:0 /R:1 /anc:1 /w:[ 31 ] /type:0
  //: joint g1380 (w71) @(526, 359) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1740 (w233) @(20, 1640) /w:[ 2 4 1 -1 ]
  //: joint g1927 (w42) @(1274, 894) /w:[ -1 2 1 4 ]
  //: joint g1454 (w219) @(416, 136) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g1287 (w215) @(337,176) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g356 (w67) @(540, 151) /anc:1 /w:[ 17 -1 18 20 ]
  //: joint g152 (w149) @(652, 143) /anc:1 /w:[ 21 -1 22 24 ]
  D_FF g1368 (.D(w76), .CP(w116), .Q(w72), .NQ(w229));   //: @(942, 2078) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>181 Ro0<9 Ro1<1 ]
  //: joint g1676 (w72) @(995, 2092) /w:[ 1 2 8 -1 ]
  //: LED g27 (w31) @(857,73) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: LED g1441 (w290) @(372,111) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g1177 (w356) @(353,274) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: joint g199 (w169) @(864, 216) /anc:1 /w:[ 7 8 10 -1 ]
  //: joint g434 (w166) @(712, 169) /anc:1 /w:[ 5 6 8 -1 ]
  //: joint g1948 (w63) @(1320, 1104) /w:[ -1 4 6 3 ]
  //: LED g636 (w181) @(715,309) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1232 (w16) @(-710, 848) /w:[ 4 42 3 -1 ]
  //: LED g1181 (w356) @(341,277) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g349 (w233) @(545, 68) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g1505 (w163) @(640,-7) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g989 (w103) @(779,134) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g2032 (w211) @(361, 1196) /w:[ 4 6 -1 3 ]
  //: joint g142 (w160) @(760, 137) /anc:1 /w:[ 35 36 -1 38 ]
  //: LED g318 (w186) @(674,351) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g829 (w0) @(484, 296) /anc:1 /w:[ 41 42 -1 44 ]
  //: comment g1977 @(742,-91)
  //: /line:"<h1 color=blue>1</h1>"
  //: /end
  //: LED g1292 (w215) @(438,186) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: joint g353 (w233) @(528, 32) /anc:1 /w:[ 31 32 -1 34 ]
  //: LED g734 (w204) @(461,297) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: LED g981 (w103) @(742,149) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: joint g1950 (w66) @(1327, 1124) /w:[ -1 6 8 5 ]
  //: joint g1871 (w34) @(-238, 1108) /w:[ 58 84 57 -1 ]
  //: joint g1449 (w219) @(364, 123) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1355 (w116) @(1127, 1995) /w:[ 120 122 119 -1 ]
  //: LED g1548 (w163) @(636,19) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g477 (w300) @(589, 430) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g937 (w211) @(362,224) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1318 (w134) @(628, 43) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g745 (w204) @(390, 330) /anc:1 /w:[ 13 14 -1 16 ]
  //: joint g1700 (w34) @(-499, 1251) /w:[ 41 42 44 -1 ]
  //: joint g299 (w286) @(782, 314) /anc:1 /w:[ 27 -1 28 30 ]
  //: joint g117 (w20) @(613, 93) /anc:1 /w:[ -1 11 12 14 ]
  //: LED g194 (w41) @(599,329) /sn:0 /R:3 /anc:1 /w:[ 7 ] /type:0
  //: LED g746 (w204) @(368,359) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g556 (w201) @(432, 432) /anc:1 /w:[ 8 10 7 -1 ]
  //: joint g767 (w296) @(504, 39) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g1733 (w34) @(-305, 1251) /w:[ 29 30 32 -1 ]
  //: joint g512 (w87) @(748, 10) /anc:1 /w:[ 15 -1 16 18 ]
  //: LED g178 (w169) @(813,204) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g426 (w32) @(579,164) /sn:0 /R:1 /anc:1 /w:[ 23 ] /type:0
  //: LED g1494 (w357) @(661,51) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: LED g1308 (w134) @(621,-20) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  D_FF g1647 (.D(w81), .CP(w116), .Q(w82), .NQ(w275));   //: @(488, 2216) /sz:(40, 56) /sn:0 /p:[ Li0>9 Li1>241 Ro0<0 Ro1<1 ]
  //: joint g1479 (w290) @(348, 93) /anc:1 /w:[ 8 10 7 -1 ]
  //: joint g1822 (w34) @(-532, 1398) /w:[ 98 97 -1 144 ]
  //: joint g1399 (w196) @(540, 456) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g456 (w28) @(610, -20) /anc:1 /w:[ 21 22 24 -1 ]
  //: LED g825 (w0) @(419,364) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1157 (w113) @(670,452) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: LED g1023 (w207) @(347,303) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g983 (w103) @(853,103) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: joint g289 (w286) @(770, 306) /anc:1 /w:[ 31 -1 32 34 ]
  //: joint g1327 (w151) @(669, 8) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1730 (w34) @(-47, 1398) /w:[ 114 128 113 -1 ]
  //: joint g1769 (w183) @(-435, 1341) /w:[ 1 2 48 -1 ]
  //: joint g412 (w27) @(513, 233) /anc:1 /w:[ 9 10 -1 12 ]
  //: LED g909 (w89) @(813,185) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g400 (w22) @(629, 291) /anc:1 /w:[ 7 8 -1 10 ]
  //: LED g389 (w166) @(688,159) /sn:0 /anc:1 /w:[ 15 ] /type:0
  //: LED g1082 (w35) @(648,467) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g310 (w186) @(654, 339) /anc:1 /w:[ 44 -1 46 43 ]
  //: LED g1704 (w36) @(251,5) /sn:0 /w:[ 1 ] /type:3
  //: joint g1966 (w93) @(1362, 1284) /w:[ -1 6 8 5 ]
  //: LED g405 (w27) @(549,230) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g1718 (w61) @(-550, 1050) /w:[ 2 4 1 -1 ]
  //: LED g605 (w265) @(419,76) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g328 (w25) @(553,292) /sn:0 /R:3 /anc:1 /w:[ 15 ] /type:0
  //: joint g976 (w103) @(842, 118) /anc:1 /w:[ 7 8 10 -1 ]
  D_FF g802 (.D(w166), .CP(w16), .Q(w19), .NQ(w94));   //: @(-566, 780) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>39 Ro0<33 Ro1<1 ]
  //: joint g1581 (w173) @(837, 261) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g394 (w22) @(638,279) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g1526 (w357) @(706, -35) /anc:1 /w:[ -1 11 12 14 ]
  //: LED g1018 (w207) @(433,267) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g820 (w0) @(440,344) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g1341 (w116) @(801, 1995) /w:[ 110 132 109 -1 ]
  //: joint g2068 (w339) @(275, 836) /w:[ 4 6 -1 3 ]
  //: joint g2061 (w169) @(295, 906) /w:[ 4 6 -1 3 ]
  //: joint g2060 (w171) @(297, 916) /w:[ 4 6 -1 3 ]
  //: LED g596 (w330) @(759,158) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g1141 (w330) @(859,129) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: LED g135 (w20) @(600,106) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g1507 (w163) @(652, -7) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1272 (w297) @(575,456) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g854 (w35) @(629,366) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g124 (w20) @(613, 130) /anc:1 /w:[ -1 23 24 26 ]
  //: joint g437 (w32) @(565, 92) /anc:1 /w:[ -1 7 8 10 ]
  //: LED g2078 (w38) @(297,5) /sn:0 /w:[ 0 ] /type:3
  //: LED g380 (w166) @(712,147) /sn:0 /anc:1 /w:[ 7 ] /type:0
  D_FF g1839 (.D(w356), .CP(w34), .Q(w283), .NQ(w370));   //: @(-36, 1481) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>181 Ro0<49 Ro1<1 ]
  D_FF g872 (.D(w11), .CP(w116), .Q(w31), .NQ(w110));   //: @(1141, 1644) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>75 Ro0<9 Ro1<1 ]
  //: LED g1600 (w174) @(822,268) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g1153 (w113) @(662,426) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: LED g284 (w317) @(506,388) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g945 (w211) @(349, 215) /anc:1 /w:[ 9 10 12 -1 ]
  //: joint g1675 (w79) @(1130, 2094) /w:[ 1 2 8 -1 ]
  //: joint g877 (w116) @(1128, 1705) /w:[ 72 74 71 -1 ]
  //: LED g1569 (w177) @(802,284) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g107 (w160) @(760,123) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g205 (w41) @(586, 280) /anc:1 /w:[ 22 24 -1 21 ]
  //: LED g707 (w332) @(799,70) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1634 (w116) @(997, 2287) /w:[ 214 224 213 -1 ]
  //: joint g661 (w202) @(485, 318) /anc:1 /w:[ 43 -1 44 46 ]
  //: joint g1926 (w132) @(1272, 884) /w:[ -1 4 6 3 ]
  //: LED g774 (w339) @(729,90) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g396 (w22) @(650,303) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g641 (w181) @(715, 321) /anc:1 /w:[ 43 -1 44 46 ]
  //: joint g2021 (w233) @(388, 1306) /w:[ 6 8 -1 5 ]
  //: LED g480 (w300) @(599,392) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: joint g1937 (w52) @(1294, 994) /w:[ -1 4 6 3 ]
  //: LED g84 (w84) @(359,37) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: joint g1598 (w173) @(862, 266) /anc:1 /w:[ -1 8 10 7 ]
  //: LED g1211 (w174) @(783,258) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g1596 (w174) @(860, 290) /anc:1 /w:[ -1 4 6 3 ]
  //: joint g723 (w298) @(769, 409) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g1448 (w352) @(388, 150) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g1669 (w69) @(800, 1942) /w:[ 6 5 8 -1 ]
  //: LED g1159 (w113) @(640,351) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g46 (w116) @(802, 1848) /w:[ 16 38 15 -1 ]
  //: LED g844 (w120) @(487,75) /sn:0 /R:1 /anc:1 /w:[ 43 ] /type:0
  //: joint g415 (w27) @(501, 238) /anc:1 /w:[ -1 8 7 26 ]
  //: joint g1304 (w134) @(631, 6) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g228 (w274) @(362, 192) /anc:1 /w:[ 13 14 16 -1 ]
  //: joint g1070 (w35) @(617, 353) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g501 (w87) @(742,-2) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g1276 (w297) @(576,443) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g1790 (w71) @(219, 1351) /w:[ 1 2 48 -1 ]
  //: joint g410 (w27) @(549, 216) /anc:1 /w:[ -1 20 19 22 ]
  //: joint g715 (w298) @(722, 356) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g1405 (w196) @(542, 443) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1158 (w113) @(662, 464) /anc:1 /w:[ 4 6 -1 3 ]
  //: joint g391 (w166) @(700, 169) /anc:1 /w:[ 9 10 -1 12 ]
  //: LED g1108 (w283) @(414,238) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g261 (w224) @(420,110) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g1929 (w40) @(1278, 914) /w:[ -1 6 8 5 ]
  //: LED g1456 (w290) @(434,135) /sn:0 /R:2 /anc:1 /w:[ 33 ] /type:0
  //: LED g1303 (w219) @(416,148) /sn:0 /R:2 /anc:1 /w:[ 33 ] /type:0
  //: LED g250 (w224) @(396,98) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g156 (w29) @(537, 189) /anc:1 /w:[ 16 -1 15 18 ]
  //: LED g701 (w332) @(740,109) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g761 (w296) @(514,75) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: joint g1350 (w116) @(998, 1995) /w:[ 116 126 115 -1 ]
  //: joint g1189 (w141) @(569, 58) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1174 (w356) @(353, 264) /anc:1 /w:[ 9 10 12 -1 ]
  //: joint g1958 (w80) @(1343, 1204) /w:[ -1 4 6 3 ]
  //: LED g16 (w41) @(599,267) /sn:0 /R:3 /anc:1 /w:[ 27 ] /type:0
  //: joint g1633 (w116) @(539, 2287) /w:[ 200 238 199 -1 ]
  //: LED g371 (w233) @(513,32) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: LED g505 (w87) @(711,46) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g1041 (w360) @(546,62) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: joint g1527 (w151) @(658, 45) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g930 (w33) @(621,455) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g788 (w339) @(729, 101) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1817 (w33) @(-112, 1346) /w:[ 1 2 48 -1 ]
  //: LED g741 (w204) @(473,289) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g308 (w186) @(698,399) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g1044 (w360) @(521,0) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g1007 (w314) @(673,397) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g553 (w201) @(474,384) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: LED g912 (w33) @(617,404) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g293 (w286) @(770,292) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1925 (w13) @(1266, 874) /w:[ -1 2 1 4 ]
  //: joint g1127 (w108) @(565, -33) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g138 (w20) @(600,118) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g188 (w169) @(764, 216) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1773 (w202) @(-377, 1489) /w:[ 1 2 48 -1 ]
  //: joint g994 (w314) @(648, 360) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g737 (w204) @(379, 338) /anc:1 /w:[ 9 10 -1 12 ]
  //: joint g1409 (w196) @(556, 367) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g498 (w87) @(757,-26) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: LED g1427 (w196) @(573,341) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: joint g672 (w202) @(474, 329) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g1542 (w357) @(697, -10) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g35 (w116) @(606, 1705) /w:[ 56 90 55 -1 ]
  //: joint g120 (w153) @(693, 59) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g1691 (w82) @(542, 2230) /w:[ 2 4 1 -1 ]
  //: joint g2062 (w89) @(293, 896) /w:[ 1 2 -1 44 ]
  //: joint g985 (w103) @(804, 134) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g226 (w274) @(388,202) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g260 (w224) @(456, 110) /anc:1 /w:[ 33 -1 34 36 ]
  //: joint g1722 (w163) @(-311, 1053) /w:[ 1 2 48 -1 ]
  //: joint g1835 (w34) @(-374, 1690) /w:[ 202 236 201 -1 ]
  D_FF g1844 (.D(w183), .CP(w34), .Q(w186), .NQ(w374));   //: @(-425, 1328) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>141 Ro0<49 Ro1<1 ]
  D_FF g1746 (.D(w35), .CP(w34), .Q(w33), .NQ(w302));   //: @(-164, 1332) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>133 Ro0<49 Ro1<1 ]
  //: joint g1584 (w174) @(759, 262) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g211 (w274) @(375, 192) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g1793 (w34) @(-176, 1108) /w:[ 60 82 59 -1 ]
  //: joint g1599 (w177) @(814, 301) /anc:1 /w:[ 19 20 22 -1 ]
  D_FF g1760 (.D(w120), .CP(w34), .Q(w296), .NQ(w321));   //: @(-102, 1625) /sz:(40, 56) /sn:0 /p:[ Li0>11 Li1>229 Ro0<0 Ro1<1 ]
  //: LED g163 (w21) @(650,233) /sn:0 /anc:1 /w:[ 31 ] /type:0
  //: LED g1296 (w215) @(349,178) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g1125 (w108) @(575,69) /sn:0 /R:1 /anc:1 /w:[ 43 ] /type:0
  //: joint g1149 (w113) @(630, 351) /anc:1 /w:[ 39 40 -1 42 ]
  D_FF g1235 (.D(w50), .CP(w116), .Q(w51), .NQ(w175));   //: @(1141, 1787) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>29 Ro0<0 Ro1<1 ]
  D_FF g1834 (.D(w33), .CP(w34), .Q(w300), .NQ(w369));   //: @(-101, 1333) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>131 Ro0<49 Ro1<1 ]
  //: joint g876 (w74) @(861, 2090) /w:[ 1 2 8 -1 ]
  //: LED g823 (w0) @(451,335) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g497 (w341) @(785,-11) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g1853 (w298) @(281, 1205) /w:[ -1 2 1 48 ]
  //: joint g1941 (w55) @(1306, 1035) /w:[ -1 4 6 3 ]
  //: joint g208 (w274) @(413, 192) /anc:1 /w:[ 29 30 32 -1 ]
  //: joint g1827 (w34) @(-239, 1398) /w:[ 108 134 107 -1 ]
  //: LED g1170 (w356) @(366,270) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: LED g262 (w224) @(360,80) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: joint g376 (w340) @(465, 258) /anc:1 /w:[ 41 42 -1 44 ]
  //: joint g1903 (w21) @(98, 648) /w:[ -1 3 4 6 ]
  //: LED g950 (w211) @(349,225) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g1006 (w314) @(648,334) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g664 (w202) @(479,340) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: LED g17 (w6) @(654,-72) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: LED g271 (w317) @(482,436) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  D_FF g1890 (.D(w304), .CP(w34), .Q(w71), .NQ(w385));   //: @(162, 1337) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>123 Ro0<49 Ro1<1 ]
  //: LED g1603 (w173) @(735,230) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: LED g572 (w204) @(485,282) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g329 (w25) @(535, 292) /anc:1 /w:[ 14 16 13 -1 ]
  //: LED g1162 (w113) @(658,413) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g716 (w298) @(760, 399) /anc:1 /w:[ 15 16 -1 18 ]
  //: LED g784 (w339) @(740,81) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: LED g270 (w317) @(500,400) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1957 (w72) @(1341, 1194) /w:[ -1 4 6 3 ]
  //: joint g358 (w233) @(540, 56) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1281 (w215) @(362, 167) /anc:1 /w:[ 13 14 16 -1 ]
  //: joint g1556 (w177) @(753, 277) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g151 (w149) @(644, 155) /anc:1 /w:[ 25 -1 26 28 ]
  //: joint g1075 (w35) @(636, 455) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g1100 (w283) @(452,231) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g1437 (w352) @(451,174) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g1485 (w352) @(375,159) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g807 (w11) @(1126, 1657) /w:[ 2 4 1 -1 ]
  //: LED g575 (w287) @(770,324) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g33 (w3) @(604, 1649) /w:[ 1 2 8 -1 ]
  //: joint g1459 (w352) @(349, 143) /anc:1 /w:[ 2 1 16 -1 ]
  //: LED g370 (w233) @(477,-40) /sn:0 /R:1 /anc:1 /w:[ 49 ] /type:0
  //: joint g1216 (w171) @(798, 235) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1122 (w108) @(551,-58) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: joint g640 (w181) @(814, 401) /anc:1 /w:[ 7 8 10 -1 ]
  assign w37 = {w32, w67, w29, w27, w25, w41, w22, w21, w19, w166, w149, w20}; //: CONCAT g1712  @(56,633) /sn:0 /R:2 /w:[ 1 33 31 31 31 31 31 27 5 0 31 31 33 ] /dr:1 /tp:1 /drp:1
  //: joint g2046 (w300) @(329, 1056) /w:[ 1 2 -1 44 ]
  //: LED g77 (w80) @(323,228) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: LED g1314 (w174) @(860,280) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: joint g1283 (w215) @(451, 176) /anc:1 /w:[ 41 42 44 -1 ]
  //: LED g342 (w186) @(686,375) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g769 (w296) @(452,-19) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g726 (w298) @(762,388) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g404 (w22) @(624, 279) /anc:1 /w:[ 12 -1 14 11 ]
  //: LED g196 (w169) @(839,204) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g566 (w181) @(803, 392) /anc:1 /w:[ 11 -1 12 14 ]
  //: LED g903 (w89) @(776,188) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1014 (w207) @(445, 252) /anc:1 /w:[ 33 34 36 -1 ]
  //: LED g246 (w224) @(456,127) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g255 (w29) @(487, 189) /anc:1 /w:[ 8 -1 7 26 ]
  D_FF g1644 (.D(w97), .CP(w116), .Q(w100), .NQ(w270));   //: @(1075, 2225) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>223 Ro0<9 Ro1<1 ]
  //: LED g1377 (w196) @(571,354) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g835 (w120) @(441, 10) /anc:1 /w:[ 17 18 -1 20 ]
  D_FF g1896 (.D(w87), .CP(w34), .Q(w341), .NQ(w387));   //: @(-35, 1044) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>79 Ro0<49 Ro1<1 ]
  //: joint g2058 (w174) @(301, 936) /w:[ 1 2 -1 44 ]
  //: LED g648 (w181) @(726,318) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g500 (w298) @(791,419) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: LED g240 (w224) @(372,86) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g652 (w181) @(726, 332) /anc:1 /w:[ 39 -1 40 42 ]
  //: LED g972 (w103) @(829,113) /sn:0 /anc:1 /w:[ 13 ] /type:0
  D_FF g1764 (.D(w89), .CP(w34), .Q(w169), .NQ(w328));   //: @(-293, 1183) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>31 Ro0<49 Ro1<1 ]
  //: joint g1970 (w97) @(1370, 1324) /w:[ -1 4 6 3 ]
  //: joint g678 (w228) @(463, 70) /anc:1 /w:[ 35 -1 36 38 ]
  //: LED g622 (w183) @(718,381) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g893 (w89) @(751,190) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g1484 (w219) @(377,138) /sn:0 /R:2 /anc:1 /w:[ 21 ] /type:0
  //: joint g1410 (w71) @(511, 395) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g298 (w286) @(806,310) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1696 (w116) @(446, 2142) /w:[ 146 145 -1 196 ]
  //: joint g1040 (w360) @(511, -49) /anc:1 /w:[ -1 7 8 10 ]
  //: joint g1715 (w32) @(1, 791) /w:[ 2 4 -1 1 ]
  //: joint g770 (w296) @(497, 27) /anc:1 /w:[ 27 28 -1 30 ]
  D_FF g1863 (.D(w215), .CP(w34), .Q(w352), .NQ(w380));   //: @(225, 1485) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>173 Ro0<11 Ro1<1 ]
  //: joint g430 (w41) @(586, 329) /anc:1 /w:[ 6 8 -1 5 ]
  //: joint g677 (w228) @(430, 42) /anc:1 /w:[ 23 -1 24 26 ]
  //: LED g614 (w265) @(467,107) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: LED g401 (w22) @(644,291) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g796 (w121) @(211, 1882) /w:[ 6 -1 8 5 ]
  //: joint g1294 (w215) @(438, 174) /anc:1 /w:[ 37 38 40 -1 ]
  //: LED g79 (w77) @(322,175) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: joint g692 (w228) @(474, 76) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g1973 (w119) @(1376, 1354) /w:[ -1 6 8 5 ]
  //: LED g1426 (w71) @(514,420) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g1046 (w360) @(551,75) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g830 (w0) @(430, 343) /anc:1 /w:[ 21 22 -1 24 ]
  //: joint g993 (w314) @(663, 397) /anc:1 /w:[ 28 30 -1 27 ]
  //: joint g1946 (w60) @(1316, 1084) /w:[ -1 4 6 3 ]
  //: joint g1709 (w19) @(-514, 794) /w:[ 30 29 32 -1 ]
  //: LED g81 (w82) @(325,122) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: joint g1180 (w356) @(429, 241) /anc:1 /w:[ 33 34 36 -1 ]
  D_FF g1729 (.D(w111), .CP(w34), .Q(w89), .NQ(w281));   //: @(-361, 1182) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>35 Ro0<49 Ro1<1 ]
  //: LED g45 (w73) @(874,283) /sn:0 /anc:1 /w:[ 3 ] /type:0
  //: LED g789 (w339) @(804,23) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g229 (w274) @(400,202) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g436 (w20) @(613, 81) /anc:1 /w:[ -1 7 8 10 ]
  PosBin60 g1974 (.pos(w45), .bin(w101));   //: @(-93, 522) /sz:(95, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: joint g1613 (w116) @(478, 2142) /w:[ 148 194 147 -1 ]
  //: joint g118 (w20) @(613, 106) /anc:1 /w:[ -1 15 16 18 ]
  //: joint g2073 (w151) @(265, 786) /w:[ 4 6 -1 3 ]
  //: LED g1455 (w219) @(403,145) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: LED g1297 (w215) @(464,189) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: comment g1987 @(615,488)
  //: /line:"<h1 color=blue>6</h1>"
  //: /end
  //: joint g1595 (w177) @(851, 313) /anc:1 /w:[ 8 -1 10 7 ]
  //: joint g1064 (w111) @(811, 174) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g478 (w300) @(599,430) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: LED g702 (w332) @(716,124) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: LED g711 (w332) @(764,94) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1172 (w356) @(441, 238) /anc:1 /w:[ 37 38 40 -1 ]
  //: joint g111 (w19) @(700, 221) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g277 (w317) @(494,412) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g11 (w5) @(600,-72) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  //: joint g1416 (w304) @(536, 377) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1383 (w71) @(520, 371) /anc:1 /w:[ 35 36 38 -1 ]
  D_FF g1856 (.D(w298), .CP(w34), .Q(w183), .NQ(w378));   //: @(-489, 1327) /sz:(40, 56) /sn:0 /p:[ Li0>49 Li1>143 Ro0<49 Ro1<1 ]
  //: joint g1351 (w116) @(931, 1995) /w:[ 114 128 113 -1 ]
  //: LED g915 (w33) @(619,429) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g1568 (w177) @(789,280) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g1414 (w304) @(530,441) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g1188 (w141) @(558, 20) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1747 (w173) @(-112, 1199) /w:[ 1 2 48 -1 ]
  //: LED g656 (w202) @(497,318) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g223 (w274) @(400, 192) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g197 (w169) @(826, 216) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g330 (w25) @(577,244) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g146 (w149) @(652,107) /sn:0 /R:1 /anc:1 /w:[ 11 ] /type:0
  //: joint g2038 (w0) @(349, 1136) /w:[ 4 6 -1 3 ]
  //: LED g452 (w28) @(600,-33) /sn:0 /R:1 /anc:1 /w:[ 19 ] /type:0
  //: joint g368 (w233) @(523, 20) /anc:1 /w:[ 27 28 -1 30 ]
  //: joint g584 (w287) @(830, 374) /anc:1 /w:[ 7 8 10 -1 ]
  D_FF g1361 (.D(w63), .CP(w116), .Q(w65), .NQ(w222));   //: @(1203, 1935) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>121 Ro0<0 Ro1<1 ]
  //: LED g417 (w32) @(573,152) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g625 (w183) @(687,333) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g227 (w274) @(450, 192) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g416 (w27) @(525, 228) /anc:1 /w:[ 13 14 -1 16 ]
  //: LED g160 (w160) @(748,129) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: joint g357 (w67) @(528, 145) /anc:1 /w:[ 13 -1 14 16 ]
  //: joint g1465 (w352) @(362, 145) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g195 (w169) @(813, 216) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g730 (w298) @(694, 323) /anc:1 /w:[ 43 44 -1 46 ]
  //: joint g1011 (w207) @(458, 247) /anc:1 /w:[ 37 38 -1 40 ]
  //: joint g1762 (w274) @(152, 1497) /w:[ 1 2 48 -1 ]
  //: LED g1266 (w219) @(440,156) /sn:0 /R:2 /anc:1 /w:[ 41 ] /type:0
  //: joint g1298 (w215) @(426, 173) /anc:1 /w:[ 33 34 36 -1 ]
  //: joint g610 (w265) @(383, 41) /anc:1 /w:[ 9 -1 10 12 ]
  //: joint g1742 (w34) @(21, 1108) /w:[ 66 76 65 -1 ]
  //: joint g1845 (w314) @(-306, 1343) /w:[ 1 2 48 -1 ]
  //: LED g14 (w3) @(628,-72) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: LED g321 (w186) @(662,327) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: joint g423 (w25) @(526, 313) /anc:1 /w:[ 6 8 -1 5 ]
  //: LED g1068 (w111) @(786,168) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g383 (w166) @(664, 186) /anc:1 /w:[ 21 22 -1 24 ]
  //: LED g1519 (w163) @(648,-46) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g362 (w233) @(537,80) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g1371 (w116) @(672, 2142) /w:[ 154 188 153 -1 ]
  //: joint g1962 (w82) @(1354, 1244) /w:[ -1 6 8 5 ]
  //: LED g1590 (w174) @(835,273) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g167 (w160) @(844,81) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g822 (w0) @(398, 371) /anc:1 /w:[ 9 10 -1 12 ]
  //: joint g906 (w89) @(776, 198) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1096 (w283) @(376, 235) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g517 (w87) @(755, -2) /anc:1 /w:[ 11 -1 12 14 ]
  //: LED g233 (w274) @(437,202) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g1565 (w174) @(835, 283) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g173 (w160) @(832, 103) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g2044 (w196) @(333, 1076) /w:[ 4 6 -1 3 ]
  //: joint g372 (w233) @(499, -28) /anc:1 /w:[ 11 12 -1 14 ]
  //: LED g759 (w296) @(460,-8) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g1358 (w116) @(866, 1995) /w:[ 112 130 111 -1 ]
  //: joint g1786 (w201) @(-437, 1488) /w:[ 1 2 48 -1 ]
  //: joint g2035 (w207) @(355, 1166) /w:[ 1 2 -1 44 ]
  //: LED g61 (w57) @(623,481) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  D_FF g1337 (.D(w47), .CP(w116), .Q(w48), .NQ(w185));   //: @(1011, 1785) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>33 Ro0<0 Ro1<1 ]
  //: joint g1801 (w34) @(-176, 1251) /w:[ 21 22 24 -1 ]
  //: LED g1204 (w141) @(563,71) /sn:0 /R:1 /anc:1 /w:[ 43 ] /type:0
  //: joint g1916 (w9) @(1250, 794) /w:[ -1 6 8 5 ]
  //: joint g1874 (w34) @(-305, 1108) /w:[ 56 86 55 -1 ]
  //: joint g1267 (w297) @(561, 468) /anc:1 /w:[ 8 10 -1 7 ]
  //: LED g441 (w340) @(465,272) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g110 (w19) @(713, 221) /anc:1 /w:[ 7 8 10 -1 ]
  //: LED g563 (w201) @(490,360) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: joint g1030 (w360) @(541, 25) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g147 (w149) @(640,131) /sn:0 /R:1 /anc:1 /w:[ 19 ] /type:0
  //: joint g1772 (w341) @(15, 1058) /w:[ 1 2 48 -1 ]
  D_FF g1843 (.D(w317), .CP(w34), .Q(w201), .NQ(w373));   //: @(-489, 1474) /sz:(40, 56) /sn:0 /p:[ Li0>49 Li1>195 Ro0<49 Ro1<1 ]
  //: joint g475 (w300) @(589, 392) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g454 (w28) @(610, 18) /anc:1 /w:[ 33 34 36 -1 ]
  //: joint g153 (w149) @(658, 131) /anc:1 /w:[ 17 -1 18 20 ]
  //: joint g1852 (w34) @(21, 1251) /w:[ 9 10 12 -1 ]
  //: joint g1219 (w16) @(-185, 848) /w:[ 20 26 19 -1 ]
  //: LED g1262 (w304) @(553,365) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g1171 (w356) @(404, 249) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g532 (w341) @(727, 77) /anc:1 /w:[ 39 -1 40 42 ]
  //: joint g1776 (w34) @(88, 1108) /w:[ 68 74 67 -1 ]
  //: LED g1207 (w141) @(548,20) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  D_FF g1622 (.D(w65), .CP(w116), .Q(w66), .NQ(w250));   //: @(489, 2071) /sz:(40, 56) /sn:0 /p:[ Li0>9 Li1>195 Ro0<0 Ro1<1 ]
  //: joint g1478 (w219) @(390, 130) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g654 (w202) @(459, 351) /anc:1 /w:[ 31 -1 32 34 ]
  //: joint g537 (w341) @(787, 0) /anc:1 /w:[ 11 -1 12 14 ]
  //: LED g69 (w68) @(407,430) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: LED g504 (w87) @(750,-14) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g573 (w287) @(782, 346) /anc:1 /w:[ 23 -1 24 26 ]
  //: joint g731 (w298) @(741, 377) /anc:1 /w:[ 23 24 -1 26 ]
  D_FF g1732 (.D(w287), .CP(w34), .Q(w181), .NQ(w288));   //: @(163, 1190) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>3 Ro0<49 Ro1<1 ]
  //: joint g1069 (w35) @(624, 391) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g1972 (w96) @(1374, 1344) /w:[ -1 4 6 3 ]
  //: joint g1920 (w10) @(1252, 804) /w:[ -1 4 6 3 ]
  //: LED g322 (w186) @(668,339) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: LED g744 (w204) @(449,304) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  D_FF g1632 (.D(w83), .CP(w116), .Q(w84), .NQ(w264));   //: @(683, 2219) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>235 Ro0<9 Ro1<1 ]
  //: joint g1254 (w171) @(862, 242) /anc:1 /w:[ -1 8 10 7 ]
  //: LED g406 (w27) @(525,242) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g743 (w204) @(473, 277) /anc:1 /w:[ 41 42 -1 44 ]
  //: joint g315 (w186) @(666, 363) /anc:1 /w:[ 35 36 -1 38 ]
  //: joint g104 (w20) @(613, 143) /anc:1 /w:[ -1 27 28 30 ]
  //: joint g1882 (w34) @(86, 1690) /w:[ 216 222 215 -1 ]
  //: LED g978 (w103) @(767,139) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: LED g133 (w20) @(600,130) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g527 (w341) @(776,0) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g627 (w183) @(675, 333) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g1446 (w352) @(388,162) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g387 (w340) @(441, 270) /anc:1 /w:[ 33 34 -1 36 ]
  //: joint g377 (w340) @(429, 275) /anc:1 /w:[ 29 30 -1 32 ]
  //: LED g961 (w64) @(587,68) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: LED g92 (w19) @(700,204) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g1396 (w71) @(532,371) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g927 (w33) @(612, 467) /anc:1 /w:[ 8 10 -1 7 ]
  //: LED g848 (w120) @(430,10) /sn:0 /R:1 /anc:1 /w:[ 19 ] /type:0
  //: LED g507 (w87) @(687,81) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1661 (w20) @(-710, 791) /w:[ 2 4 1 -1 ]
  //: LED g1589 (w174) @(848,276) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g170 (w160) @(808, 113) /anc:1 /w:[ 19 20 -1 22 ]
  //: LED g618 (w183) @(695,345) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g66 (w63) @(495,471) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g12 (w34) @(-532, 1108) /w:[ 48 94 -1 47 ]
  //: LED g543 (w120) @(448,32) /sn:0 /R:1 /anc:1 /w:[ 27 ] /type:0
  D_FF g1767 (.D(w103), .CP(w34), .Q(w330), .NQ(w334));   //: @(-488, 1180) /sz:(40, 56) /sn:0 /p:[ Li0>49 Li1>43 Ro0<49 Ro1<1 ]
  //: joint g1662 (w5) @(540, 1591) /w:[ -1 4 10 3 ]
  //: LED g108 (w160) @(772,117) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1200 (w141) @(562, 33) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g134 (w20) @(600,93) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g326 (w25) @(571,256) /sn:0 /R:3 /anc:1 /w:[ 27 ] /type:0
  //: LED g1413 (w304) @(527,454) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g2033 (w283) @(359, 1186) /w:[ 4 6 -1 3 ]
  //: joint g552 (w201) @(476, 360) /anc:1 /w:[ 31 -1 32 34 ]
  D_FF g1812 (.D(w233), .CP(w34), .Q(w360), .NQ(w361));   //: @(31, 1627) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>225 Ro0<49 Ro1<1 ]
  //: joint g996 (w314) @(684, 447) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g1798 (w34) @(-48, 1690) /w:[ 212 226 211 -1 ]
  D_FF g1230 (.D(w20), .CP(w16), .Q(w149), .NQ(w145));   //: @(-697, 778) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>43 Ro0<33 Ro1<1 ]
  //: LED g1145 (w330) @(796,147) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g773 (w339) @(783, 55) /anc:1 /w:[ 19 20 -1 22 ]
  //: joint g1666 (w53) @(604, 1939) /w:[ 1 2 8 -1 ]
  //: joint g335 (w25) @(541, 280) /anc:1 /w:[ 18 20 17 -1 ]
  //: joint g1547 (w357) @(692, 2) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1058 (w111) @(850,156) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g793 (w116) @(673, 1848) /w:[ 12 42 11 -1 ]
  //: LED g225 (w274) @(425,202) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g1673 (w60) @(1065, 1946) /w:[ 1 2 8 -1 ]
  //: joint g440 (w27) @(489, 238) /anc:1 /w:[ 6 -1 5 28 ]
  //: LED g177 (w169) @(751,204) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: LED g192 (w169) @(788,204) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1334 (w304) @(517, 454) /anc:1 /w:[ 7 8 10 -1 ]
  //: LED g901 (w89) @(738,191) /sn:0 /anc:1 /w:[ 43 ] /type:0
  //: LED g1551 (w177) @(753,265) /sn:0 /anc:1 /w:[ 41 ] /type:0
  D_FF g1340 (.D(w46), .CP(w116), .Q(w73), .NQ(w191));   //: @(878, 1783) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>37 Ro0<9 Ro1<1 ]
  //: joint g1911 (w19) @(96, 658) /w:[ -1 2 1 28 ]
  //: LED g312 (w186) @(716,435) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: joint g653 (w202) @(414, 406) /anc:1 /w:[ 11 -1 12 14 ]
  //: LED g286 (w286) @(818,316) /sn:0 /anc:1 /w:[ 17 ] /type:0
  D_FF g1752 (.D(w296), .CP(w34), .Q(w233), .NQ(w313));   //: @(-37, 1626) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>227 Ro0<0 Ro1<1 ]
  //: LED g683 (w228) @(452,72) /sn:0 /R:2 /anc:1 /w:[ 33 ] /type:0
  //: LED g25 (w11) @(845,36) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g466 (w28) @(600,30) /sn:0 /R:1 /anc:1 /w:[ 39 ] /type:0
  //: LED g1552 (w174) @(733,243) /sn:0 /anc:1 /w:[ 43 ] /type:0
  D_FF g1808 (.D(w201), .CP(w34), .Q(w202), .NQ(w359));   //: @(-425, 1475) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>193 Ro0<49 Ro1<1 ]
  //: joint g1275 (w297) @(567, 417) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g100 (w41) @(586, 267) /anc:1 /w:[ 26 28 -1 25 ]
  //: joint g942 (w211) @(375, 213) /anc:1 /w:[ 17 18 20 -1 ]
  //: joint g2042 (w71) @(337, 1096) /w:[ 4 6 -1 3 ]
  //: joint g253 (w224) @(384, 74) /anc:1 /w:[ 12 11 -1 42 ]
  //: LED g1385 (w196) @(565,379) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: joint g1476 (w219) @(428, 139) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g155 (w149) @(669, 107) /anc:1 /w:[ 9 -1 10 12 ]
  //: joint g123 (w153) @(729, -13) /anc:1 /w:[ 15 -1 16 18 ]
  //: LED g1106 (w283) @(401,240) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: LED g1486 (w290) @(385,117) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: LED g1290 (w163) @(651,-58) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: LED g1265 (w297) @(579,417) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1758 (w151) @(-239, 1054) /w:[ 1 2 48 -1 ]
  //: LED g243 (w29) @(475,202) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: joint g1618 (w116) @(739, 2142) /w:[ 156 186 155 -1 ]
  //: joint g1964 (w83) @(1358, 1264) /w:[ -1 4 6 3 ]
  //: LED g355 (w67) @(528,163) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1238 (w171) @(850, 240) /anc:1 /w:[ 11 12 14 -1 ]
  D_FF g1763 (.D(w357), .CP(w34), .Q(w153), .NQ(w327));   //: @(-163, 1042) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>83 Ro0<49 Ro1<1 ]
  //: LED g987 (w103) @(792,129) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g1060 (w111) @(748,175) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g828 (w0) @(408,373) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g252 (w224) @(420, 94) /anc:1 /w:[ 21 -1 22 24 ]
  //: joint g1554 (w177) @(827, 305) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1541 (w163) @(662, -58) /anc:1 /w:[ -1 7 8 10 ]
  //: joint g1898 (w34) @(-500, 1545) /w:[ 148 194 147 -1 ]
  //: LED g623 (w183) @(741,416) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g99 (w153) @(701, 35) /anc:1 /w:[ 31 -1 32 34 ]
  D_FF g1714 (.D(w290), .CP(w34), .Q(w224), .NQ(w269));   //: @(-363, 1621) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>237 Ro0<49 Ro1<1 ]
  //: LED g951 (w64) @(577,-58) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: LED g1029 (w207) @(421,272) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: joint g1194 (w141) @(539, -43) /anc:1 /w:[ 8 7 -1 10 ]
  //: joint g1930 (w44) @(1280, 924) /w:[ -1 6 8 5 ]
  //: joint g2031 (w274) @(363, 1206) /w:[ 4 6 -1 3 ]
  //: comment g1980 @(237,-45) /sn:0
  //: /line:"<h1 color=red>HH:MM:SS</h1>"
  //: /end
  //: LED g103 (w149) @(628,155) /sn:0 /R:1 /anc:1 /w:[ 27 ] /type:0
  //: joint g1829 (w34) @(-46, 1108) /w:[ 64 78 63 -1 ]
  //: joint g10 (w116) @(479, 1705) /w:[ 52 94 51 -1 ]
  //: joint g1771 (w34) @(150, 1108) /w:[ 70 72 69 -1 ]
  //: joint g1079 (w35) @(637, 467) /anc:1 /w:[ 8 10 -1 7 ]
  //: LED g1558 (w173) @(761,235) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: joint g1672 (w59) @(998, 1945) /w:[ 1 2 8 -1 ]
  D_FF g1847 (.D(w297), .CP(w34), .Q(w196), .NQ(w376));   //: @(32, 1335) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>127 Ro0<49 Ro1<1 ]
  //: joint g1615 (w116) @(1193, 2142) /w:[ 170 172 169 -1 ]
  //: GROUND g9 (w4) @(388,1722) /sn:0 /R:1 /w:[ 0 ]
  D_FF g1620 (.D(w77), .CP(w116), .Q(w81), .NQ(w247));   //: @(1203, 2082) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>173 Ro0<0 Ro1<1 ]
  //: joint g898 (w89) @(764, 199) /anc:1 /w:[ 35 36 38 -1 ]
  D_FF g1749 (.D(w174), .CP(w34), .Q(w177), .NQ(w307));   //: @(-35, 1187) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>15 Ro0<49 Ro1<1 ]
  //: joint g660 (w202) @(405, 417) /anc:1 /w:[ 8 10 7 -1 ]
  //: joint g1686 (w90) @(927, 2236) /w:[ 2 4 1 -1 ]
  //: LED g474 (w300) @(599,342) /sn:0 /R:3 /anc:1 /w:[ 43 ] /type:0
  //: joint g2070 (w87) @(271, 816) /w:[ 1 2 -1 44 ]
  //: LED g42 (w44) @(876,230) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: LED g1442 (w352) @(438,171) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g1067 (w111) @(837, 168) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g862 (w108) @(570,43) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g1027 (w207) @(408,277) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: comment g1985 @(863,345)
  //: /line:"<h1 color=blue>4</h1>"
  //: /end
  //: joint g1728 (w207) @(-117, 1493) /w:[ 46 45 48 -1 ]
  //: LED g612 (w265) @(478,116) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g435 (w149) @(675, 95) /anc:1 /w:[ -1 5 6 8 ]
  //: LED g22 (w24) @(795,-23) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: LED g70 (w70) @(376,404) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: joint g651 (w181) @(781, 376) /anc:1 /w:[ 19 -1 20 22 ]
  //: LED g114 (w153) @(682,47) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g378 (w340) @(369,320) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  D_FF g879 (.D(w14), .CP(w116), .Q(w24), .NQ(w123));   //: @(943, 1641) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>81 Ro0<9 Ro1<1 ]
  //: joint g164 (w21) @(662, 257) /anc:1 /w:[ -1 26 28 25 ]
  //: LED g165 (w160) @(784,111) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g1373 (w304) @(523,466) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  D_FF g1641 (.D(w86), .CP(w116), .Q(w83), .NQ(w268));   //: @(615, 2218) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>237 Ro0<9 Ro1<1 ]
  //: joint g496 (w341) @(796, -11) /anc:1 /w:[ -1 7 8 10 ]
  //: joint g140 (w153) @(740, -37) /anc:1 /w:[ -1 7 8 10 ]
  //: LED g1533 (w151) @(669,-31) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g1870 (w296) @(-51, 1639) /w:[ 2 4 1 -1 ]
  //: joint g1594 (w174) @(809, 276) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g1534 (w163) @(638,6) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  D_FF g1621 (.D(w72), .CP(w116), .Q(w80), .NQ(w248));   //: @(1010, 2079) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>179 Ro0<9 Ro1<1 ]
  //: joint g706 (w332) @(787, 94) /anc:1 /w:[ 23 24 -1 26 ]
  //: joint g1240 (w171) @(748, 230) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1183 (w356) @(392, 252) /anc:1 /w:[ 21 22 24 -1 ]
  //: joint g1420 (w304) @(513, 466) /anc:1 /w:[ 4 6 -1 3 ]
  D_FF g1331 (.D(w42), .CP(w116), .Q(w156), .NQ(w176));   //: @(617, 1779) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>45 Ro0<9 Ro1<1 ]
  //: joint g1838 (w34) @(87, 1398) /w:[ 118 124 117 -1 ]
  //: joint g1854 (w34) @(150, 1251) /w:[ 1 2 4 -1 ]
  //: joint g965 (w64) @(588, -46) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g590 (w287) @(734,301) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: LED g130 (w153) @(699,11) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g1311 (w134) @(626,-58) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: frame g1976 @(-545,1011) /sn:0 /wi:860 /ht:700 /tx:"sequence of flip-flops as shift register"
  D_FF g1825 (.D(w330), .CP(w34), .Q(w111), .NQ(w366));   //: @(-424, 1181) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>39 Ro0<49 Ro1<1 ]
  //: LED g1268 (w297) @(583,367) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  PosBin12 g1913 (.pos(w37), .bin(w36));   //: @(-93, 568) /sz:(100, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: LED g1165 (w113) @(655,401) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: frame g1994 @(223,-96) /sn:0 /wi:161 /ht:121 /tx:"Digital clock"
  //: LED g1085 (w35) @(624,340) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g1400 (w196) @(551,456) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g230 (w41) @(599,317) /sn:0 /R:3 /anc:1 /w:[ 11 ] /type:0
  D_FF g1781 (.D(w61), .CP(w34), .Q(w28), .NQ(w345));   //: @(-488, 1037) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>93 Ro0<53 Ro1<1 ]
  //: joint g1935 (w50) @(1290, 974) /w:[ -1 6 8 5 ]
  //: joint g753 (w296) @(482, 4) /anc:1 /w:[ 19 20 -1 22 ]
  D_FF g1645 (.D(w96), .CP(w116), .Q(w119), .NQ(w135));   //: @(1202, 2227) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>219 Ro0<0 Ro1<1 ]
  //: LED g1054 (w111) @(824,161) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g1309 (w134) @(617,31) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g1094 (w283) @(376,245) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1021 (w207) @(458,257) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: joint g2069 (w341) @(273, 826) /w:[ 4 6 -1 3 ]
  //: LED g762 (w296) @(467,4) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g1091 (w283) @(363,248) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g870 (w116) @(1066, 1705) /w:[ 70 76 69 -1 ]
  //: joint g1654 (w44) @(803, 1795) /w:[ 2 4 1 -1 ]
  //: LED g297 (w286) @(746,281) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: joint g320 (w186) @(695, 423) /anc:1 /w:[ 15 16 -1 18 ]
  //: LED g1393 (w71) @(519,408) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g1857 (w297) @(20, 1348) /w:[ 1 2 48 -1 ]
  //: joint g1884 (w34) @(-111, 1251) /w:[ 17 18 20 -1 ]
  //: joint g2019 (w141) @(392, 1326) /w:[ 1 2 -1 44 ]
  //: LED g23 (w12) @(826,4) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: joint g1787 (w211) @(84, 1496) /w:[ 1 2 48 -1 ]
  //: frame g2000 @(334,1849) /sn:0 /wi:101 /ht:40 /tx:"Start Stop AND"
  //: LED g470 (w28) @(600,5) /sn:0 /R:1 /anc:1 /w:[ 31 ] /type:0
  //: joint g1037 (w360) @(526, -12) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g1184 (w356) @(467,240) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g1451 (w352) @(401, 152) /anc:1 /w:[ 29 30 32 -1 ]
  //: joint g973 (w103) @(792, 139) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1253 (w171) @(811, 236) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1136 (w330) @(771,155) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: joint g671 (w202) @(430, 384) /anc:1 /w:[ 19 -1 20 22 ]
  //: LED g1500 (w357) @(691,-23) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g399 (w340) @(453,278) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: LED g136 (w153) @(723,-37) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: LED g591 (w287) @(758,316) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: LED g190 (w169) @(764,204) /sn:0 /anc:1 /w:[ 41 ] /type:0
  //: joint g1951 (w68) @(1329, 1134) /w:[ -1 4 6 3 ]
  //: joint g1225 (w16) @(-449, 848) /w:[ 12 34 11 -1 ]
  //: LED g1137 (w330) @(847,132) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g2047 (w33) @(327, 1046) /w:[ 4 6 -1 3 ]
  //: joint g502 (w87) @(725, 46) /anc:1 /w:[ 27 -1 28 30 ]
  //: joint g1432 (w219) @(351, 120) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g1610 (w116) @(931, 2142) /w:[ 162 180 161 -1 ]
  //: joint g1968 (w90) @(1366, 1304) /w:[ -1 6 8 5 ]
  //: LED g781 (w339) @(718,100) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1567 (w173) @(798, 254) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1024 (w207) @(396,282) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1490 (w290) @(471,150) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g1270 (w297) @(571, 367) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g2017 (w64) @(396, 1346) /w:[ 4 6 -1 3 ]
  //: joint g1329 (w304) @(530, 402) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g96 (w116) @(1066, 1848) /w:[ 24 30 23 -1 ]
  //: joint g1367 (w116) @(1065, 2142) /w:[ 166 176 165 -1 ]
  //: joint g1636 (w116) @(604, 2287) /w:[ 202 236 201 -1 ]
  //: LED g812 (w0) @(484,306) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g1461 (w290) @(458, 133) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1084 (w35) @(628, 416) /anc:1 /w:[ 23 24 26 -1 ]
  D_FF g808 (.D(w31), .CP(w116), .Q(w13), .NQ(w106));   //: @(1204, 1645) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>73 Ro0<7 Ro1<1 ]
  //: LED g171 (w21) @(638,227) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g586 (w287) @(818, 367) /anc:1 /w:[ 11 -1 12 14 ]
  //: joint g1101 (w283) @(427, 225) /anc:1 /w:[ 33 34 36 -1 ]
  D_FF g1799 (.D(w196), .CP(w34), .Q(w304), .NQ(w353));   //: @(98, 1336) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>125 Ro0<49 Ro1<1 ]
  //: joint g1820 (w34) @(149, 1545) /w:[ 168 174 167 -1 ]
  //: joint g1509 (w151) @(676, -18) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g1697 (w16) @(-772, 848) /w:[ 2 44 1 -1 ]
  //: joint g1789 (w290) @(-376, 1634) /w:[ 1 2 48 -1 ]
  //: joint g398 (w22) @(612, 255) /anc:1 /w:[ 20 -1 22 19 ]
  //: LED g360 (w233) @(525,56) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g463 (w28) @(610, 30) /anc:1 /w:[ 37 38 40 -1 ]
  //: joint g43 (w116) @(740, 1705) /w:[ 60 86 59 -1 ]
  //: LED g587 (w287) @(806,347) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g361 (w233) @(504, -16) /anc:1 /w:[ 15 16 -1 18 ]
  //: joint g1346 (w116) @(672, 1995) /w:[ 106 136 105 -1 ]
  //: joint g1354 (w116) @(478, 1995) /w:[ 100 142 99 -1 ]
  //: joint g1813 (w287) @(152, 1203) /w:[ 1 2 48 -1 ]
  //: joint g2063 (w111) @(291, 886) /w:[ 1 2 -1 44 ]
  //: joint g1169 (w356) @(454, 234) /anc:1 /w:[ 41 42 -1 44 ]
  //: joint g2075 (w134) @(261, 766) /w:[ 4 6 -1 3 ]
  //: LED g513 (w87) @(703,58) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g2022 (w296) @(386, 1296) /w:[ 6 8 -1 5 ]
  //: LED g941 (w211) @(463,216) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: LED g975 (w103) @(816,119) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: joint g1559 (w177) @(765, 283) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1566 (w174) @(822, 280) /anc:1 /w:[ 15 16 18 -1 ]
  //: comment g1983 @(327,-63) /sn:0
  //: /line:"<h3 color=blue>RUN</h3>"
  //: /end
  //: LED g1606 (w177) @(728,256) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: joint g1901 (w20) @(90, 688) /w:[ -1 6 32 5 ]
  //: joint g698 (w332) @(740, 120) /anc:1 /w:[ 39 40 -1 42 ]
  //: LED g214 (w41) @(599,292) /sn:0 /R:3 /anc:1 /w:[ 19 ] /type:0
  //: LED g1545 (w357) @(685,-10) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: LED g933 (w211) @(450,217) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g1072 (w35) @(626, 404) /anc:1 /w:[ 28 30 -1 27 ]
  //: LED g471 (w28) @(600,42) /sn:0 /R:1 /anc:1 /w:[ 43 ] /type:0
  //: LED g859 (w356) @(441,248) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: joint g1438 (w290) @(372, 101) /anc:1 /w:[ 16 -1 15 46 ]
  D_FF g1754 (.D(w173), .CP(w34), .Q(w174), .NQ(w315));   //: @(-100, 1186) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>19 Ro0<49 Ro1<1 ]
  //: joint g606 (w265) @(478, 102) /anc:1 /w:[ 42 41 -1 44 ]
  //: LED g1032 (w360) @(510,-25) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g154 (w149) @(664, 119) /anc:1 /w:[ 13 -1 14 16 ]
  //: LED g530 (w341) @(722,66) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g1150 (w113) @(666,439) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g418 (w32) @(561,128) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: joint g750 (w204) @(425, 306) /anc:1 /w:[ 25 26 -1 28 ]
  //: joint g1942 (w69) @(1308, 1044) /w:[ -1 1 2 4 ]
  //: frame g1996 @(-156,454) /sn:0 /wi:191 /ht:173 /tx:" position to binary conversion"
  //: joint g1899 (w67) @(-59, 801) /w:[ 1 2 32 -1 ]
  //: LED g1392 (w71) @(523,395) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g1190 (w141) @(533,-30) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: LED g354 (w233) @(483,-28) /sn:0 /R:1 /anc:1 /w:[ 13 ] /type:0
  //: joint g907 (w89) @(864, 191) /anc:1 /w:[ -1 4 6 3 ]
  //: joint g1423 (w71) @(502, 420) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g76 (w72) @(324,255) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: joint g841 (w120) @(423, -10) /anc:1 /w:[ 3 4 14 -1 ]
  //: LED g647 (w181) @(781,363) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g1132 (w330) @(759, 168) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g1430 (w71) @(547,334) /sn:0 /R:3 /anc:1 /w:[ 47 ] /type:0
  //: LED g364 (w233) @(519,44) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g1944 (w58) @(1312, 1064) /w:[ -1 4 6 3 ]
  //: LED g998 (w314) @(663,372) /sn:0 /R:3 /anc:1 /w:[ 37 ] /type:0
  //: LED g687 (w228) @(419,45) /sn:0 /R:2 /anc:1 /w:[ 21 ] /type:0
  //: joint g1954 (w75) @(1335, 1164) /w:[ -1 6 8 5 ]
  //: joint g631 (w183) @(697, 369) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g359 (w233) @(533, 44) /anc:1 /w:[ 35 36 -1 38 ]
  //: LED g929 (w33) @(618,416) /sn:0 /R:3 /anc:1 /w:[ 25 ] /type:0
  //: joint g468 (w28) @(610, 55) /anc:1 /w:[ 45 46 48 -1 ]
  D_FF g801 (.D(w6), .CP(w116), .Q(w9), .NQ(w92));   //: @(685, 1637) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>89 Ro0<0 Ro1<1 ]
  //: joint g1291 (w215) @(337, 164) /anc:1 /w:[ 8 -1 7 46 ]
  //: LED g1489 (w352) @(414,166) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g1564 (w173) @(811, 256) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1963 (w86) @(1356, 1254) /w:[ -1 4 6 3 ]
  _GGOR2 #(6) g6 (.I0(w7), .I1(w119), .Z(w114));   //: @(271,1812) /sn:0 /R:1 /w:[ 7 3 0 ]
  //: joint g882 (w16) @(-252, 848) /w:[ 18 28 17 -1 ]
  //: joint g922 (w33) @(609, 429) /anc:1 /w:[ 19 20 22 -1 ]
  D_FF g1357 (.D(w53), .CP(w116), .Q(w56), .NQ(w218));   //: @(616, 1926) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>139 Ro0<9 Ro1<1 ]
  //: joint g980 (w103) @(853, 114) /anc:1 /w:[ 3 4 6 -1 ]
  //: joint g1510 (w163) @(650, 6) /anc:1 /w:[ 27 28 30 -1 ]
  D_FF g1627 (.D(w90), .CP(w116), .Q(w95), .NQ(w254));   //: @(941, 2223) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>227 Ro0<0 Ro1<1 ]
  //: LED g149 (w160) @(724,141) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: joint g2037 (w204) @(351, 1146) /w:[ 4 6 -1 3 ]
  //: joint g338 (w67) @(552, 159) /anc:1 /w:[ 22 21 -1 24 ]
  //: LED g1103 (w283) @(389,242) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g1185 (w356) @(404,259) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  D_FF g1879 (.D(w300), .CP(w34), .Q(w297), .NQ(w382));   //: @(-36, 1334) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>129 Ro0<49 Ro1<1 ]
  //: LED g48 (w47) @(865,309) /sn:0 /anc:1 /w:[ 7 ] /type:0
  //: joint g1959 (w79) @(1345, 1214) /w:[ -1 4 6 3 ]
  //: joint g1836 (w34) @(87, 1545) /w:[ 166 176 165 -1 ]
  //: LED g1580 (w177) @(741,261) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1218 (w16) @(-123, 848) /w:[ 22 24 21 -1 ]
  //: joint g300 (w286) @(818, 334) /anc:1 /w:[ 15 -1 16 18 ]
  //: joint g1131 (w330) @(796, 157) /anc:1 /w:[ 27 28 30 -1 ]
  _GGOR2 #(6) g1698 (.I0(w18), .I1(w4), .Z(w23));   //: @(408,1685) /sn:0 /w:[ 0 1 0 ]
  //: LED g560 (w201) @(514,325) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: LED g581 (w287) @(782,332) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g232 (w29) @(537,202) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1324 (w134) @(623,-33) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  D_FF g1619 (.D(w80), .CP(w116), .Q(w79), .NQ(w245));   //: @(1076, 2080) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>177 Ro0<9 Ro1<1 ]
  //: joint g1953 (w193) @(1333, 1154) /w:[ -1 1 2 4 ]
  //: joint g1575 (w173) @(850, 263) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g41 (w116) @(802, 1705) /w:[ 62 84 61 -1 ]
  //: joint g1692 (w84) @(736, 2233) /w:[ 1 2 8 -1 ]
  //: joint g1753 (w169) @(-240, 1197) /w:[ 1 2 48 -1 ]
  //: LED g1328 (w304) @(545,389) /sn:0 /R:3 /anc:1 /w:[ 29 ] /type:0
  //: LED g90 (w97) @(495,-63) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  D_FF g1805 (.D(w28), .CP(w34), .Q(w134), .NQ(w358));   //: @(-424, 1038) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>91 Ro0<49 Ro1<1 ]
  //: joint g1864 (w34) @(-240, 1690) /w:[ 206 232 205 -1 ]
  //: LED g924 (w33) @(616,391) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g1381 (w71) @(508,433) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  D_FF g1646 (.D(w95), .CP(w116), .Q(w97), .NQ(w273));   //: @(1009, 2224) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>225 Ro0<9 Ro1<1 ]
  //: joint g1872 (w34) @(149, 1398) /w:[ 120 122 119 -1 ]
  //: joint g1694 (w116) @(446, 1848) /w:[ 4 50 -1 3 ]
  //: joint g1516 (w163) @(655, -20) /anc:1 /w:[ 19 20 22 -1 ]
  //: joint g1135 (w330) @(821, 150) /anc:1 /w:[ 19 20 22 -1 ]
  D_FF g1217 (.D(w44), .CP(w116), .Q(w46), .NQ(w170));   //: @(815, 1782) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>39 Ro0<0 Ro1<1 ]
  //: joint g1922 (w11) @(1262, 854) /w:[ -1 6 8 5 ]
  signal g1330 (.p(w7), .p1(w17), .p2(w8), .fdbks(fdbk60), .clk(w121));   //: @(67, 1856) /sz:(129, 107) /sn:0 /p:[ Lo0<0 Lo1<1 Lo2<0 Ro0<17 Ro1<9 ]
  //: LED g148 (w160) @(796,105) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: joint g461 (w28) @(610, -7) /anc:1 /w:[ 25 26 28 -1 ]
  //: LED g1549 (w357) @(652,76) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g1814 (w34) @(-532, 1251) /w:[ 45 46 -1 96 ]
  //: joint g1850 (w34) @(20, 1545) /w:[ 164 178 163 -1 ]
  //: LED g943 (w211) @(425,219) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: joint g926 (w33) @(605, 379) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g467 (w28) @(600,-7) /sn:0 /R:1 /anc:1 /w:[ 27 ] /type:0
  //: LED g1433 (w219) @(339,126) /sn:0 /R:2 /anc:1 /w:[ 49 ] /type:0
  //: joint g1688 (w93) @(802, 2234) /w:[ 2 4 1 -1 ]
  //: LED g189 (w169) @(738,204) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: LED g995 (w314) @(683,421) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  D_FF g1344 (.D(w55), .CP(w116), .Q(w69), .NQ(w206));   //: @(750, 1928) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>135 Ro0<9 Ro1<1 ]
  //: LED g212 (w274) @(375,202) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g1313 (w134) @(620,-7) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g509 (w87) @(696,70) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: joint g309 (w186) @(704, 447) /anc:1 /w:[ 8 -1 10 7 ]
  //: LED g1057 (w111) @(773,171) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1518 (w163) @(659, -46) /anc:1 /w:[ -1 11 12 14 ]
  //: LED g742 (w204) @(402,336) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g539 (w341) @(767,11) /sn:0 /R:1 /anc:1 /w:[ 17 ] /type:0
  //: LED g595 (w339) @(707,109) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: joint g403 (w22) @(634, 303) /anc:1 /w:[ 4 -1 6 3 ]
  //: LED g1597 (w177) @(777,275) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1785 (w153) @(-113, 1056) /w:[ 1 2 48 -1 ]
  //: LED g534 (w341) @(704,88) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: joint g977 (w103) @(816, 129) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g409 (w27) @(537,236) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: LED g295 (w286) @(734,275) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g851 (w193) @(735, 2088) /w:[ 6 5 8 -1 ]
  //: joint g1022 (w207) @(433, 257) /anc:1 /w:[ 29 30 32 -1 ]
  //: LED g643 (w181) @(748,336) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g2051 (w186) @(319, 1006) /w:[ 4 6 -1 3 ]
  //: LED g846 (w120) @(478,64) /sn:0 /R:1 /anc:1 /w:[ 39 ] /type:0
  //: LED g73 (w19) @(650,204) /sn:0 /anc:1 /w:[ 27 ] /type:0
  //: joint g327 (w186) @(683, 399) /anc:1 /w:[ 23 24 -1 26 ]
  //: LED g928 (w33) @(614,367) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g1586 (w177) @(789, 292) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g74 (w74) @(333,308) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: LED g421 (w32) @(567,140) /sn:0 /R:1 /anc:1 /w:[ 27 ] /type:0
  //: LED g36 (w42) @(876,150) /sn:0 /anc:1 /w:[ 3 ] /type:0
  //: LED g216 (w274) @(349,202) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g1123 (w108) @(561,-7) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g1191 (w141) @(554, 8) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1851 (w34) @(-439, 1690) /w:[ 200 238 199 -1 ]
  //: LED g144 (w149) @(646,119) /sn:0 /R:1 /anc:1 /w:[ 15 ] /type:0
  //: joint g1195 (w141) @(547, -17) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1332 (w116) @(867, 1848) /w:[ 18 36 17 -1 ]
  D_FF g853 (.D(w22), .CP(w16), .Q(w41), .NQ(w105));   //: @(-373, 783) /sz:(40, 56) /sn:0 /p:[ Li0>31 Li1>33 Ro0<33 Ro1<1 ]
  //: LED g1147 (w330) @(784,151) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: joint g1585 (w173) @(761, 247) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g528 (w341) @(695,98) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g708 (w332) @(776, 100) /anc:1 /w:[ 27 28 -1 30 ]
  //: joint g1339 (w13) @(1259, 1659) /w:[ -1 5 6 8 ]
  //: LED g1142 (w330) @(808,144) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g382 (w166) @(676,165) /sn:0 /anc:1 /w:[ 19 ] /type:0
  //: joint g525 (w341) @(761, 33) /anc:1 /w:[ 23 -1 24 26 ]
  //: joint g1682 (w100) @(1126, 2239) /w:[ 1 2 8 -1 ]
  _GGMUX2 #(8, 8) g13 (.I0(w17), .I1(w2), .S(fdbk60), .Z(w61));   //: @(-616,1050) /sn:0 /R:1 /w:[ 0 1 0 0 ] /ss:0 /do:0
  //: LED g55 (w54) @(765,451) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g1280 (w215) @(401, 171) /anc:1 /w:[ 25 26 28 -1 ]
  //: joint g604 (w265) @(443, 78) /anc:1 /w:[ 29 -1 30 32 ]
  //: joint g905 (w89) @(852, 192) /anc:1 /w:[ 7 8 10 -1 ]
  //: LED g1205 (w141) @(544,8) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: joint g176 (w160) @(844, 99) /anc:1 /w:[ 7 8 -1 10 ]
  //: joint g637 (w181) @(770, 366) /anc:1 /w:[ 23 -1 24 26 ]
  //: joint g1717 (w28) @(-438, 1003) /w:[ -1 4 50 3 ]
  //: comment g1992 @(459,-92)
  //: /line:"<h1 color=blue>11</h1>"
  //: /end
  //: joint g1 (w6) @(667, 1650) /w:[ 1 2 8 -1 ]
  //: LED g344 (w233) @(507,20) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: joint g550 (w201) @(469, 372) /anc:1 /w:[ 27 -1 28 30 ]
  //: LED g992 (w314) @(689,434) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: joint g2054 (w181) @(309, 976) /w:[ 4 6 -1 3 ]
  //: LED g1602 (w177) @(814,289) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: LED g1117 (w108) @(568,31) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g1095 (w283) @(350, 240) /anc:1 /w:[ 9 10 12 -1 ]
  //: joint g1140 (w330) @(771, 165) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g306 (w286) @(842,328) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: LED g1531 (w357) @(700,-47) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: LED g132 (w153) @(687,35) /sn:0 /R:1 /anc:1 /w:[ 33 ] /type:0
  //: joint g113 (w19) @(676, 221) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g414 (w27) @(561,224) /sn:0 /R:2 /anc:1 /w:[ 21 ] /type:0
  //: LED g1012 (w207) @(371,293) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: LED g1458 (w219) @(428,151) /sn:0 /R:2 /anc:1 /w:[ 37 ] /type:0
  //: joint g1684 (w95) @(998, 2237) /w:[ 2 4 1 -1 ]
  //: comment g1991 @(313,56)
  //: /line:"<h1 color=blue>10</h1>"
  //: /end
  //: joint g1325 (w134) @(636, -46) /anc:1 /w:[ -1 11 12 14 ]
  //: joint g1099 (w283) @(338, 241) /anc:1 /w:[ 8 -1 7 46 ]
  D_FF g1748 (.D(w71), .CP(w34), .Q(w317), .NQ(w306));   //: @(225, 1338) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>121 Ro0<0 Ro1<1 ]
  D_FF g1369 (.D(w193), .CP(w116), .Q(w75), .NQ(w232));   //: @(750, 2075) /sz:(40, 56) /sn:0 /p:[ Li0>7 Li1>187 Ro0<0 Ro1<1 ]
  //: LED g31 (w132) @(873,124) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: LED g20 (w15) @(730,-51) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: joint g169 (w160) @(820, 108) /anc:1 /w:[ 15 16 -1 18 ]
  //: LED g869 (w89) @(864,181) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: joint g967 (w64) @(587, -58) /anc:1 /w:[ -1 7 8 10 ]
  //: LED g68 (w66) @(436,445) /sn:0 /R:3 /anc:1 /w:[ 7 ] /type:0
  //: LED g772 (w339) @(751,71) /sn:0 /anc:1 /w:[ 33 ] /type:0
  D_FF g795 (.D(w10), .CP(w116), .Q(w15), .NQ(w85));   //: @(815, 1639) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>85 Ro0<9 Ro1<1 ]
  //: LED g694 (w332) @(787,78) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: LED g703 (w332) @(728,117) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: LED g544 (w296) @(521,87) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: joint g179 (w169) @(776, 216) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g52 (w19) @(676,204) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: LED g838 (w120) @(506,97) /sn:0 /R:1 /anc:1 /w:[ 49 ] /type:0
  //: LED g1001 (w314) @(653,347) /sn:0 /R:3 /anc:1 /w:[ 45 ] /type:0
  //: joint g1830 (w339) @(84, 1059) /w:[ 1 2 48 -1 ]
  //: LED g704 (w332) @(752,102) /sn:0 /anc:1 /w:[ 37 ] /type:0
  D_FF g1228 (.D(w149), .CP(w16), .Q(w166), .NQ(w143));   //: @(-634, 779) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>41 Ro0<33 Ro1<1 ]
  //: LED g1197 (w141) @(530,-43) /sn:0 /R:1 /anc:1 /w:[ 9 ] /type:0
  //: joint g1611 (w116) @(605, 2142) /w:[ 152 190 151 -1 ]
  //: joint g47 (w15) @(865, 1653) /w:[ 1 2 8 -1 ]
  //: joint g1146 (w330) @(834, 146) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1658 (w66) @(541, 2085) /w:[ 2 4 1 -1 ]
  //: joint g105 (w160) @(784, 127) /anc:1 /w:[ 27 28 -1 30 ]
  //: LED g247 (w29) @(500,202) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: joint g988 (w103) @(829, 123) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g1828 (w34) @(20, 1398) /w:[ 116 126 115 -1 ]
  //: LED g710 (w332) @(833,47) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g918 (w33) @(604, 367) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g311 (w186) @(671, 375) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g116 (w20) @(613, 118) /anc:1 /w:[ -1 19 20 22 ]
  //: joint g990 (w314) @(658, 384) /anc:1 /w:[ 32 34 -1 31 ]
  //: LED g1512 (w357) @(680,2) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: joint g337 (w186) @(690, 411) /anc:1 /w:[ 19 20 -1 22 ]
  //: joint g278 (w317) @(490, 388) /anc:1 /w:[ 28 30 27 -1 ]
  //: joint g439 (w29) @(475, 189) /anc:1 /w:[ 6 -1 5 28 ]
  //: LED g697 (w332) @(822,55) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g1469 (w352) @(438, 159) /anc:1 /w:[ 41 42 44 -1 ]
  //: joint g224 (w41) @(586, 292) /anc:1 /w:[ 18 20 -1 17 ]
  //: LED g892 (w89) @(801,186) /sn:0 /anc:1 /w:[ 25 ] /type:0
  //: comment g1993 @(587,-111)
  //: /line:"<h1 color=blue>12</h1>"
  //: /end
  //: LED g449 (w340) @(429,290) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: LED g910 (w89) @(852,182) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g1467 (w290) @(360, 96) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g331 (w186) @(704,411) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g220 (w41) @(599,280) /sn:0 /R:3 /anc:1 /w:[ 23 ] /type:0
  D_FF g1842 (.D(w360), .CP(w34), .Q(w141), .NQ(w372));   //: @(97, 1628) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>223 Ro0<49 Ro1<1 ]
  //: joint g1113 (w108) @(580, 43) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1033 (w360) @(536, 12) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g679 (w228) @(441, 52) /anc:1 /w:[ 27 -1 28 30 ]
  //: LED g931 (w211) @(337,226) /sn:0 /R:2 /anc:1 /w:[ 47 ] /type:0
  //: LED g569 (w202) @(416,417) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1401 (w71) @(530, 347) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g1129 (w330) @(746, 172) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g98 (w153) @(664,83) /sn:0 /R:1 /anc:1 /w:[ 47 ] /type:0
  //: LED g944 (w211) @(413,220) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: joint g880 (w12) @(1062, 1656) /w:[ 1 2 8 -1 ]
  //: LED g317 (w25) @(541,316) /sn:0 /R:3 /anc:1 /w:[ 7 ] /type:0
  //: joint g775 (w339) @(740, 92) /anc:1 /w:[ 35 36 -1 38 ]
  //: LED g425 (w32) @(555,116) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: LED g87 (w91) @(399,-22) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  //: LED g78 (w79) @(322,202) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: LED g1263 (w297) @(573,468) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1529 (w357) @(688, 15) /anc:1 /w:[ 27 28 30 -1 ]
  //: LED g1074 (w35) @(641,429) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: LED g1063 (w111) @(811,164) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g258 (w29) @(512, 189) /anc:1 /w:[ 12 -1 11 22 ]
  //: LED g1605 (w173) @(785,240) /sn:0 /anc:1 /w:[ 33 ] /type:0
  //: LED g143 (w149) @(634,143) /sn:0 /R:1 /anc:1 /w:[ 23 ] /type:0
  //: joint g765 (w296) @(473, -8) /anc:1 /w:[ 15 16 -1 18 ]
  //: joint g162 (w21) @(674, 264) /anc:1 /w:[ -1 22 24 21 ]
  //: joint g791 (w339) @(814, 26) /anc:1 /w:[ 7 8 -1 10 ]
  //: joint g127 (w153) @(717, 11) /anc:1 /w:[ 23 -1 24 26 ]
  //: LED g633 (w183) @(749,427) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0
  //: LED g443 (w340) @(381,314) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: LED g367 (w233) @(495,-4) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g958 (w64) @(595, 42) /anc:1 /w:[ 39 40 42 -1 ]
  //: joint g1723 (w186) @(-374, 1342) /w:[ 1 2 48 -1 ]
  //: LED g62 (w58) @(599,482) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: LED g1161 (w113) @(673,464) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: LED g63 (w59) @(570,483) /sn:0 /R:3 /anc:1 /w:[ 5 ] /type:0
  //: joint g1317 (w134) @(630, 19) /anc:1 /w:[ 31 32 34 -1 ]
  //: joint g695 (w332) @(728, 129) /anc:1 /w:[ 43 44 -1 46 ]
  //: LED g1445 (w352) @(426,168) /sn:0 /R:2 /anc:1 /w:[ 39 ] /type:0
  //: LED g234 (w224) @(384,92) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: joint g175 (w160) @(796, 120) /anc:1 /w:[ 23 24 -1 26 ]
  //: LED g574 (w287) @(746,308) /sn:0 /anc:1 /w:[ 37 ] /type:0
  //: LED g588 (w287) @(723,292) /sn:0 /anc:1 /w:[ 45 ] /type:0
  //: joint g1702 (fdbk60) @(-616, 1090) /w:[ -1 1 2 8 ]
  //: LED g85 (w93) @(375,7) /sn:0 /R:2 /anc:1 /w:[ 7 ] /type:0
  //: joint g1450 (w219) @(377, 126) /anc:1 /w:[ 19 20 22 -1 ]
  //: LED g385 (w166) @(664,171) /sn:0 /anc:1 /w:[ 23 ] /type:0
  //: frame g1999 @(-10,1825) /sn:0 /wi:240 /ht:175 /tx:"Signal generator"
  //: LED g589 (w287) @(830,362) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: LED g1462 (w219) @(390,142) /sn:0 /R:2 /anc:1 /w:[ 25 ] /type:0
  //: joint g1389 (w304) @(520, 441) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g313 (w186) @(659, 351) /anc:1 /w:[ 39 40 -1 42 ]
  //: LED g101 (w27) @(489,260) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: LED g384 (w166) @(700,153) /sn:0 /anc:1 /w:[ 11 ] /type:0
  //: LED g1199 (w141) @(559,58) /sn:0 /R:1 /anc:1 /w:[ 41 ] /type:0
  //: joint g1434 (w219) @(453, 148) /anc:1 /w:[ 43 44 46 -1 ]
  //: joint g432 (w21) @(710, 276) /anc:1 /w:[ 2 1 12 -1 ]
  //: joint g235 (w224) @(360, 63) /anc:1 /w:[ 8 -1 7 46 ]
  //: joint g184 (w21) @(698, 274) /anc:1 /w:[ 13 14 16 -1 ]
  //: joint g1931 (w46) @(1282, 934) /w:[ -1 6 8 5 ]
  //: joint g1322 (w134) @(629, 31) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g219 (w274) @(425, 192) /anc:1 /w:[ 33 34 36 -1 ]
  //: LED g479 (w300) @(599,355) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g920 (w33) @(610, 442) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g237 (w224) @(432, 102) /anc:1 /w:[ 25 -1 26 28 ]
  //: joint g186 (w21) @(650, 249) /anc:1 /w:[ -1 30 32 29 ]
  //: joint g533 (w341) @(771, 22) /anc:1 /w:[ 19 -1 20 22 ]
  //: joint g1961 (w81) @(1349, 1234) /w:[ -1 4 6 3 ]
  //: joint g2076 (w28) @(259, 756) /w:[ 6 8 -1 5 ]
  //: joint g1411 (w196) @(559, 354) /anc:1 /w:[ 43 44 46 -1 ]
  //: LED g429 (w340) @(477,266) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: joint g268 (w317) @(498, 376) /anc:1 /w:[ 32 34 31 -1 ]
  //: LED g1062 (w111) @(862,154) /sn:0 /anc:1 /w:[ 5 ] /type:0
  //: LED g292 (w286) @(830,322) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: joint g438 (w67) @(492, 128) /anc:1 /w:[ 6 -1 5 28 ]
  //: joint g1391 (w196) @(549, 404) /anc:1 /w:[ 27 28 30 -1 ]
  //: joint g1048 (w360) @(520, -25) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g787 (w339) @(751, 82) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g1876 (w34) @(-306, 1398) /w:[ 106 136 105 -1 ]
  //: joint g1909 (w27) @(106, 608) /w:[ -1 4 30 3 ]
  //: joint g121 (w160) @(772, 132) /anc:1 /w:[ 31 32 -1 34 ]
  //: joint g1005 (w314) @(668, 409) /anc:1 /w:[ 24 26 -1 23 ]
  //: joint g1774 (w34) @(-307, 1690) /w:[ 204 234 203 -1 ]
  //: LED g1435 (w290) @(446,141) /sn:0 /R:2 /anc:1 /w:[ 37 ] /type:0
  //: joint g712 (w332) @(822, 68) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g1222 (w116) @(932, 1848) /w:[ 20 34 19 -1 ]
  //: LED g1286 (w352) @(337,151) /sn:0 /R:2 /anc:1 /w:[ 15 ] /type:0
  //: joint g1152 (w113) @(634, 364) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g392 (w166) @(676, 179) /anc:1 /w:[ 17 18 -1 20 ]
  D_FF g1336 (.D(w51), .CP(w116), .Q(w52), .NQ(w184));   //: @(1204, 1788) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>27 Ro0<9 Ro1<1 ]
  //: joint g7 (w7) @(291, 1854) /w:[ -1 4 6 3 ]
  //: joint g343 (w186) @(700, 435) /anc:1 /w:[ 11 12 -1 14 ]
  //: joint g603 (w265) @(395, 48) /anc:1 /w:[ 13 -1 14 16 ]
  //: joint g1107 (w283) @(363, 238) /anc:1 /w:[ 13 14 16 -1 ]
  //: LED g778 (w339) @(762,62) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: joint g1653 (w40) @(738, 1794) /w:[ 2 4 1 -1 ]
  //: joint g1869 (w113) @(-241, 1344) /w:[ 46 45 48 -1 ]
  //: LED g729 (w298) @(771,399) /sn:0 /R:3 /anc:1 /w:[ 17 ] /type:0
  //: LED g986 (w103) @(729,154) /sn:0 /anc:1 /w:[ 43 ] /type:0
  D_FF g1624 (.D(w74), .CP(w116), .Q(w76), .NQ(w251));   //: @(877, 2077) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>183 Ro0<9 Ro1<1 ]
  //: joint g1800 (w265) @(-242, 1636) /w:[ 1 2 48 -1 ]
  //: joint g1356 (w77) @(1191, 2095) /w:[ 2 4 1 -1 ]
  //: joint g1390 (w304) @(523, 428) /anc:1 /w:[ 15 16 18 -1 ]
  //: LED g83 (w83) @(346,74) /sn:0 /R:2 /anc:1 /w:[ 5 ] /type:0
  //: joint g273 (w317) @(500, 364) /anc:1 /w:[ 36 38 -1 35 ]
  //: joint g1659 (w68) @(601, 2086) /w:[ 1 2 8 -1 ]
  //: joint g2043 (w304) @(335, 1086) /w:[ 1 2 -1 44 ]
  //: comment g1988 @(448,464)
  //: /line:"<h1 color=blue>7</h1>"
  //: /end
  D_FF g809 (.D(w24), .CP(w116), .Q(w12), .NQ(w107));   //: @(1011, 1642) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>79 Ro0<9 Ro1<1 ]
  //: LED g668 (w202) @(488,329) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: LED g740 (w204) @(414,328) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g856 (w314) @(658,360) /sn:0 /R:3 /anc:1 /w:[ 41 ] /type:0
  //: joint g248 (w29) @(525, 189) /anc:1 /w:[ 14 -1 13 20 ]
  //: joint g814 (w0) @(451, 324) /anc:1 /w:[ 29 30 -1 32 ]
  //: joint g1683 (w96) @(1190, 2240) /w:[ 1 2 8 -1 ]
  //: joint g1689 (w83) @(670, 2232) /w:[ 1 2 8 -1 ]
  //: LED g159 (w149) @(658,95) /sn:0 /R:1 /anc:1 /w:[ 7 ] /type:0
  //: joint g1826 (w34) @(-437, 1251) /w:[ 37 38 40 -1 ]
  //: comment g1981 @(238,-63) /sn:0
  //: /line:"<h3 color=blue>+1 h</h3>"
  //: /end
  //: joint g1034 (w360) @(551, 49) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g571 (w0) @(430,355) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: joint g1877 (w111) @(-370, 1195) /w:[ 46 45 48 -1 ]
  //: LED g645 (w181) @(792,372) /sn:0 /anc:1 /w:[ 17 ] /type:0
  //: LED g1576 (w173) @(850,252) /sn:0 /anc:1 /w:[ 13 ] /type:0
  //: LED g1035 (w360) @(516,-12) /sn:0 /R:1 /anc:1 /w:[ 21 ] /type:0
  //: joint g490 (w300) @(589, 443) /anc:1 /w:[ 11 12 14 -1 ]
  //: LED g339 (w67) @(492,145) /sn:0 /R:2 /anc:1 /w:[ 29 ] /type:0
  //: LED g826 (w0) @(462,325) /sn:0 /R:2 /anc:1 /w:[ 35 ] /type:0
  //: LED g979 (w103) @(842,108) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g2057 (w177) @(303, 946) /w:[ 4 6 -1 3 ]
  //: joint g1912 (w149) @(92, 678) /w:[ -1 4 30 3 ]
  //: joint g1307 (w134) @(626, 56) /anc:1 /w:[ -1 43 44 46 ]
  //: LED g1133 (w330) @(821,140) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: LED g1421 (w71) @(528,383) /sn:0 /R:3 /anc:1 /w:[ 33 ] /type:0
  //: LED g128 (w153) @(693,23) /sn:0 /R:1 /anc:1 /w:[ 29 ] /type:0
  //: joint g954 (w64) @(591, -7) /anc:1 /w:[ 23 24 26 -1 ]
  //: joint g1192 (w141) @(565, 45) /anc:1 /w:[ 35 36 38 -1 ]
  //: LED g158 (w21) @(674,245) /sn:0 /anc:1 /w:[ 23 ] /type:0
  //: joint g1387 (w196) @(553, 379) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g600 (w265) @(407, 55) /anc:1 /w:[ 17 -1 18 20 ]
  D_FF g1794 (.D(w141), .CP(w34), .Q(w108), .NQ(w350));   //: @(161, 1629) /sz:(40, 56) /sn:0 /p:[ Li0>47 Li1>221 Ro0<49 Ro1<1 ]
  //: joint g1915 (w3) @(1246, 774) /w:[ -1 4 6 3 ]
  D_FF g884 (.D(w19), .CP(w16), .Q(w21), .NQ(w78));   //: @(-500, 781) /sz:(40, 56) /sn:0 /p:[ Li0>31 Li1>37 Ro0<11 Ro1<1 ]
  //: joint g1407 (w71) @(493, 445) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g699 (w332) @(752, 113) /anc:1 /w:[ 35 36 -1 38 ]
  //: joint g947 (w211) @(337, 216) /anc:1 /w:[ 8 -1 7 46 ]
  //: joint g161 (w160) @(736, 149) /anc:1 /w:[ 43 44 -1 46 ]
  //: joint g934 (w211) @(388, 212) /anc:1 /w:[ 21 22 24 -1 ]
  //: joint g1491 (w151) @(682, -44) /anc:1 /w:[ -1 11 12 14 ]
  //: LED g445 (w340) @(393,308) /sn:0 /R:2 /anc:1 /w:[ 19 ] /type:0
  //: LED g363 (w233) @(531,68) /sn:0 /R:1 /anc:1 /w:[ 45 ] /type:0
  //: LED g764 (w296) @(499,51) /sn:0 /R:1 /anc:1 /w:[ 37 ] /type:0
  //: LED g1477 (w219) @(453,160) /sn:0 /R:2 /anc:1 /w:[ 45 ] /type:0
  //: LED g1003 (w314) @(699,458) /sn:0 /R:3 /anc:1 /w:[ 9 ] /type:0
  //: joint g1020 (w207) @(347, 292) /anc:1 /w:[ 4 -1 3 42 ]
  //: joint g1887 (w34) @(-373, 1398) /w:[ 104 138 103 -1 ]
  //: joint g32 (w31) @(1192, 1658) /w:[ 1 2 8 -1 ]
  //: joint g1073 (w35) @(619, 366) /anc:1 /w:[ 39 40 42 -1 ]
  //: LED g408 (w27) @(501,254) /sn:0 /R:2 /anc:1 /w:[ 27 ] /type:0
  //: LED g1201 (w141) @(526,-55) /sn:0 /R:1 /anc:1 /w:[ 5 ] /type:0
  //: joint g1237 (w116) @(1128, 1848) /w:[ 26 28 25 -1 ]
  D_FF g1363 (.D(w52), .CP(w116), .Q(w54), .NQ(w225));   //: @(489, 1924) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>143 Ro0<9 Ro1<1 ]
  //: joint g1674 (w62) @(1131, 1947) /w:[ 1 2 8 -1 ]
  //: LED g1210 (w173) @(862,255) /sn:0 /anc:1 /w:[ 9 ] /type:0
  //: joint g1388 (w196) @(547, 417) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g1126 (w108) @(563,5) /sn:0 /R:1 /anc:1 /w:[ 25 ] /type:0
  //: LED g615 (w265) @(443,92) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: joint g790 (w339) @(762, 73) /anc:1 /w:[ 27 28 -1 30 ]
  //: joint g718 (w298) @(731, 367) /anc:1 /w:[ 27 28 -1 30 ]
  //: joint g959 (w64) @(593, 18) /anc:1 /w:[ 31 32 34 -1 ]
  //: LED g71 (w193) @(355,368) /sn:0 /R:2 /anc:1 /w:[ 0 ] /type:0
  //: LED g1591 (w173) @(798,242) /sn:0 /anc:1 /w:[ 29 ] /type:0
  //: LED g749 (w204) @(379,351) /sn:0 /R:2 /anc:1 /w:[ 11 ] /type:0
  //: joint g1008 (w314) @(679, 434) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1408 (w304) @(541, 365) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1002 (w314) @(653, 372) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g1053 (w111) @(761, 183) /anc:1 /w:[ 35 36 38 -1 ]
  //: joint g748 (w204) @(461, 286) /anc:1 /w:[ 37 38 -1 40 ]
  //: joint g1932 (w73) @(1284, 944) /w:[ -1 2 1 4 ]
  //: joint g1888 (w34) @(-372, 1108) /w:[ 54 88 53 -1 ]
  assign w45 = {w119, w96, w100, w97, w95, w90, w91, w93, w84, w83, w86, w82, w81, w77, w79, w80, w72, w76, w74, w75, w193, w70, w68, w66, w65, w63, w62, w60, w59, w58, w57, w69, w55, w56, w53, w54, w52, w51, w50, w48, w47, w73, w46, w44, w40, w156, w42, w132, w13, w31, w11, w12, w24, w14, w15, w10, w9, w6, w3, w5}; //: CONCAT g1713  @(1192,1059) /sn:0 /R:2 /w:[ 1 9 7 7 7 9 9 9 9 7 7 7 9 7 9 7 7 7 7 7 9 3 9 7 9 7 7 7 7 7 7 7 3 7 7 7 7 7 9 9 9 9 0 9 9 9 0 0 7 0 7 9 7 7 0 7 7 9 7 7 9 ] /dr:0 /tp:0 /drp:1
  D_FF g1859 (.D(w151), .CP(w34), .Q(w357), .NQ(w379));   //: @(-227, 1041) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>85 Ro0<49 Ro1<1 ]
  //: LED g1241 (w171) @(735,217) /sn:0 /anc:1 /w:[ 47 ] /type:0
  //: LED g949 (w211) @(388,222) /sn:0 /R:2 /anc:1 /w:[ 23 ] /type:0
  //: LED g1179 (w356) @(454,244) /sn:0 /R:2 /anc:1 /w:[ 43 ] /type:0
  //: LED g782 (w339) @(783,42) /sn:0 /anc:1 /w:[ 21 ] /type:0
  //: joint g971 (w103) @(742, 159) /anc:1 /w:[ 39 40 -1 42 ]
  //: joint g1705 (fdbk60) @(-837, 893) /w:[ -1 4 6 3 ]
  //: joint g489 (w300) @(589, 355) /anc:1 /w:[ 39 40 42 -1 ]
  D_FF g1832 (.D(w153), .CP(w34), .Q(w87), .NQ(w368));   //: @(-100, 1043) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>81 Ro0<49 Ro1<1 ]
  _GGAND2 #(6) g1707 (.I0(w61), .I1(w28), .Z(w30));   //: @(-547,981) /sn:0 /R:1 /w:[ 5 51 1 ]
  //: joint g1154 (w113) @(660, 452) /anc:1 /w:[ 7 8 10 -1 ]
  //: LED g667 (w202) @(443,384) /sn:0 /R:3 /anc:1 /w:[ 21 ] /type:0
  //: joint g551 (w201) @(446, 408) /anc:1 /w:[ 15 -1 16 18 ]
  //: LED g1475 (w352) @(401,164) /sn:0 /R:2 /anc:1 /w:[ 31 ] /type:0
  //: joint g1703 (w149) @(-646, 792) /w:[ 1 2 32 -1 ]
  //: joint g1846 (w34) @(-499, 1108) /w:[ 50 92 49 -1 ]
  //: joint g2029 (w352) @(367, 1226) /w:[ 6 5 -1 8 ]
  D_FF g1725 (.D(w283), .CP(w34), .Q(w211), .NQ(w277));   //: @(32, 1482) /sz:(40, 56) /sn:0 /p:[ Li0>0 Li1>179 Ro0<49 Ro1<1 ]
  //: joint g2027 (w290) @(376, 1246) /w:[ 4 6 -1 3 ]
  //: joint g209 (w274) @(337, 192) /anc:1 /w:[ 8 -1 7 46 ]
  //: joint g2064 (w330) @(289, 876) /w:[ 4 6 -1 3 ]
  //: joint g1087 (w35) @(634, 442) /anc:1 /w:[ 15 16 18 -1 ]
  //: joint g1891 (w219) @(-436, 1633) /w:[ 2 4 1 -1 ]
  D_FF g1720 (.D(w219), .CP(w34), .Q(w290), .NQ(w261));   //: @(-426, 1620) /sz:(40, 56) /sn:0 /p:[ Li0>3 Li1>239 Ro0<49 Ro1<1 ]
  //: joint g1583 (w177) @(839, 310) /anc:1 /w:[ 11 12 14 -1 ]
  //: joint g486 (w300) @(589, 405) /anc:1 /w:[ 23 24 26 -1 ]
  //: LED g728 (w298) @(781,409) /sn:0 /R:3 /anc:1 /w:[ 13 ] /type:0

endmodule
//: /netlistEnd

//: /netlistBegin NorMos
module NorMos(B, A, Z);
//: interface  /sz:(60, 40) /bd:[ Ri0>B(16/40) Ri1>A(28/40) Lo0<Z(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(144,182)(210,182){1}
//: {2}(214,182)(260,182){3}
//: {4}(212,184)(212,235)(227,235){5}
supply1 w114;    //: /sn:0 {0}(274,126)(274,113){1}
input A;    //: /sn:0 {0}(150,134)(247,134){1}
//: {2}(251,134)(260,134){3}
//: {4}(249,136)(249,236)(299,236){5}
output Z;    //: /sn:0 {0}(313,228)(313,213){1}
//: {2}(315,211)(390,211)(390,211)(405,211){3}
//: {4}(313,209)(313,208)(276,208){5}
//: {6}(274,206)(274,191){7}
//: {8}(272,208)(241,208)(241,227){9}
supply0 w116;    //: /sn:0 {0}(313,245)(313,261)(276,261){1}
//: {2}(272,261)(241,261)(241,244){3}
//: {4}(274,263)(274,272){5}
wire w121;    //: /sn:0 {0}(274,143)(274,174){1}
//: enddecls

  //: IN g3 (B) @(142,182) /sn:0 /w:[ 0 ]
  //: joint g1987 (w116) @(274, 261) /w:[ 1 -1 2 4 ]
  //: joint g1989 (A) @(249, 134) /w:[ 2 -1 1 4 ]
  //: IN g2 (A) @(148,134) /sn:0 /w:[ 0 ]
  //: joint g1992 (Z) @(274, 208) /w:[ 5 6 8 -1 ]
  _GGPMOS #(2, 1) g1995 (.Z(Z), .S(w121), .G(B));   //: @(268,182) /sn:0 /w:[ 7 1 3 ]
  //: OUT g1 (Z) @(402,211) /sn:0 /w:[ 3 ]
  //: VDD g1982 (w114) @(285,113) /sn:0 /w:[ 1 ]
  //: GROUND g1988 (w116) @(274,278) /sn:0 /w:[ 5 ]
  //: joint g1985 (B) @(212, 182) /w:[ 2 -1 1 4 ]
  _GGNMOS #(2, 1) g1983 (.Z(Z), .S(w116), .G(A));   //: @(307,236) /sn:0 /w:[ 0 0 5 ]
  _GGNMOS #(2, 1) g1990 (.Z(Z), .S(w116), .G(B));   //: @(235,235) /sn:0 /w:[ 9 3 5 ]
  //: joint g0 (Z) @(313, 211) /w:[ 2 4 -1 1 ]
  _GGPMOS #(2, 1) g1993 (.Z(w121), .S(w114), .G(A));   //: @(268,134) /sn:0 /w:[ 0 0 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin PosBin60
module PosBin60(pos, bin);
//: interface  /sz:(95, 40) /bd:[ Li0>pos[59:0](18/40) Ro0<bin[5:0](16/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [5:0] bin;    //: /sn:0 {0}(3370,475)(3266,475)(3266,475)(#:3243,475){1}
input [59:0] pos;    //: /sn:0 {0}(#:-25,452)(-2,452)(-2,452)(#:19,452){1}
wire w32;    //: /sn:0 {0}(532,262)(511,262)(511,262)(491,262){1}
wire w160;    //: /sn:0 {0}(1672,385)(1630,385)(1630,385)(1642,385){1}
wire w73;    //: /sn:0 {0}(639,244)(692,244)(692,249)(706,249){1}
wire w96;    //: /sn:0 {0}(25,737)(3089,737)(3089,512){1}
//: {2}(3091,510)(3101,510)(3101,510)(3114,510){3}
//: {4}(3089,508)(3089,498)(3089,498)(3089,498){5}
//: {6}(3091,496)(3101,496)(3101,496)(3114,496){7}
//: {8}(3089,494)(3089,484){9}
//: {10}(3091,482)(3114,482){11}
//: {12}(3089,480)(3089,473)(3089,473)(3089,460)(3089,460)(3089,454)(3104,454)(3104,454)(3114,454){13}
wire w45;    //: /sn:0 {0}(490,220)(510,220)(510,225)(609,225){1}
wire w244;    //: /sn:0 {0}(2968,434)(2996,434)(2996,444)(3114,444){1}
wire w166;    //: /sn:0 {0}(3144,505)(3142,505)(3142,505)(3177,505){1}
wire w134;    //: /sn:0 {0}(1248,314)(1089,314)(1089,306)(991,306)(991,293)(987,293){1}
wire w141;    //: /sn:0 {0}(639,271)(686,271)(686,286)(818,286)(818,299)(908,299)(908,308)(1016,308){1}
wire w220;    //: /sn:0 {0}(2723,470)(2710,470)(2710,470)(2754,470){1}
wire w14;    //: /sn:0 {0}(188,218)(164,218)(164,218)(200,218){1}
wire w218;    //: /sn:0 {0}(2693,409)(2658,409)(2658,409)(2672,409){1}
wire w16;    //: /sn:0 {0}(231,195)(241,195){1}
wire w56;    //: /sn:0 {0}(1177,346)(1166,346)(1166,346)(1155,346){1}
//: {2}(1153,344)(1153,340)(1153,340)(1153,335){3}
//: {4}(1155,333)(1166,333)(1166,333)(1177,333){5}
//: {6}(1153,331)(1153,321)(1153,321)(1153,311){7}
//: {8}(1155,309)(1172,309)(1172,309)(1177,309){9}
//: {10}(1153,307)(1153,295)(1177,295){11}
//: {12}(1153,348)(1153,427)(25,427){13}
wire w179;    //: /sn:0 {0}(2122,392)(2087,392)(2087,392)(2090,392){1}
wire w4;    //: /sn:0 {0}(85,188)(155,188)(155,199)(158,199){1}
wire w19;    //: /sn:0 {0}(656,286)(635,286)(635,317)(25,317){1}
wire w81;    //: /sn:0 {0}(25,627)(2436,627)(2436,457){1}
//: {2}(2438,455)(2448,455)(2448,455)(2461,455){3}
//: {4}(2436,453)(2436,443)(2436,443)(2436,429){5}
//: {6}(2438,427)(2461,427){7}
//: {8}(2436,425)(2436,418)(2436,418)(2436,415){9}
//: {10}(2438,413)(2449,413)(2449,413)(2461,413){11}
//: {12}(2436,411)(2436,405)(2436,405)(2436,401){13}
//: {14}(2438,399)(2451,399)(2451,399)(2461,399){15}
//: {16}(2436,397)(2436,385)(2461,385){17}
wire w89;    //: /sn:0 {0}(987,263)(997,263)(997,271)(1056,271)(1056,278)(1070,278){1}
wire w195;    //: /sn:0 {0}(2243,402)(2238,402)(2238,402)(2277,402){1}
wire w38;    //: /sn:0 {0}(25,257)(270,257)(270,254){1}
//: {2}(272,252)(277,252)(277,252)(286,252){3}
//: {4}(270,250)(270,224)(288,224){5}
wire w182;    //: /sn:0 {0}(2243,374)(2255,374)(2255,384)(2401,384){1}
wire w180;    //: /sn:0 {0}(2243,430)(2238,430)(2238,430)(2277,430){1}
wire w152;    //: /sn:0 {0}(1456,316)(1439,316)(1439,316)(1422,316){1}
wire w183;    //: /sn:0 {0}(2090,350)(2185,350)(2185,355)(2213,355){1}
wire w3;    //: /sn:0 {0}(25,247)(227,247)(227,249){1}
//: {2}(229,247)(231,247)(231,247)(239,247){3}
//: {4}(227,245)(227,205)(241,205){5}
wire w181;    //: /sn:0 {0}(3177,449)(3142,449)(3142,449)(3144,449){1}
wire w151;    //: /sn:0 {0}(1207,304)(1260,304)(1260,311)(1392,311){1}
wire w0;    //: /sn:0 {0}(231,209)(259,209)(259,214)(288,214){1}
wire w127;    //: /sn:0 {0}(1248,328)(1227,328)(1227,328)(1207,328){1}
wire w233;    //: /sn:0 {0}(2938,485)(2889,485)(2889,485)(2908,485){1}
wire w133;    //: /sn:0 {0}(25,437)(1223,437)(1223,353){1}
//: {2}(1225,351)(1236,351)(1236,351)(1248,351){3}
//: {4}(1223,349)(1223,345)(1223,345)(1223,340){5}
//: {6}(1225,338)(1236,338)(1236,338)(1248,338){7}
//: {8}(1223,336)(1223,324)(1248,324){9}
wire w171;    //: /sn:0 {0}(1872,358)(1823,358)(1823,358)(1835,358){1}
wire w168;    //: /sn:0 {0}(1578,310)(1622,310)(1622,315)(1672,315){1}
wire w111;    //: /sn:0 {0}(1456,300)(1368,300)(1368,295)(1347,295){1}
wire w104;    //: /sn:0 {0}(873,253)(935,253)(935,258)(957,258){1}
wire w204;    //: /sn:0 {0}(2523,450)(2474,450)(2474,450)(2491,450){1}
wire w75;    //: /sn:0 {0}(25,557)(1967,557)(1967,422){1}
//: {2}(1969,420)(1980,420)(1980,420)(1990,420){3}
//: {4}(1967,418)(1967,392)(1990,392){5}
wire w237;    //: /sn:0 {0}(2784,461)(2785,461)(2785,461)(2817,461){1}
wire w54;    //: /sn:0 {0}(25,397)(998,397)(998,333){1}
//: {2}(1000,331)(1016,331){3}
//: {4}(998,329)(998,318)(1016,318){5}
wire w209;    //: /sn:0 {0}(2642,404)(2590,404)(2590,394)(2491,394){1}
wire w67;    //: /sn:0 {0}(25,337)(693,337)(693,303){1}
//: {2}(695,301)(697,301)(697,301)(705,301){3}
//: {4}(693,299)(693,259)(706,259){5}
wire w215;    //: /sn:0 {0}(2491,422)(2513,422)(2513,506)(2958,506)(2958,462)(2987,462){1}
wire w90;    //: /sn:0 {0}(25,697)(2853,697)(2853,492){1}
//: {2}(2855,490)(2865,490)(2865,490)(2878,490){3}
//: {4}(2853,488)(2853,478)(2853,478)(2853,478){5}
//: {6}(2855,476)(2865,476)(2865,476)(2878,476){7}
//: {8}(2853,474)(2853,453)(2853,453)(2853,450){9}
//: {10}(2855,448)(2866,448)(2866,448)(2878,448){11}
//: {12}(2853,446)(2853,440)(2853,440)(2853,434)(2868,434)(2868,434)(2878,434){13}
wire w176;    //: /sn:0 {0}(3144,491)(3142,491)(3142,491)(3177,491){1}
wire w156;    //: /sn:0 {0}(532,272)(523,272)(523,272)(515,272){1}
//: {2}(513,270)(513,270)(513,270)(513,260){3}
//: {4}(515,258)(522,258)(522,258)(532,258){5}
//: {6}(513,256)(513,244)(532,244){7}
//: {8}(513,274)(513,275)(498,275)(498,297)(25,297){9}
wire w167;    //: /sn:0 {0}(1760,353)(1753,353)(1753,353)(1805,353){1}
wire w41;    //: /sn:0 {0}(25,747)(3152,747)(3152,517){1}
//: {2}(3154,515)(3164,515)(3164,515)(3177,515){3}
//: {4}(3152,513)(3152,503)(3152,503)(3152,503){5}
//: {6}(3154,501)(3164,501)(3164,501)(3177,501){7}
//: {8}(3152,499)(3152,489){9}
//: {10}(3154,487)(3177,487){11}
//: {12}(3152,485)(3152,478)(3152,478)(3152,465)(3152,465)(3152,461){13}
//: {14}(3154,459)(3167,459)(3167,459)(3177,459){15}
//: {16}(3152,457)(3152,445)(3177,445){17}
wire w36;    //: /sn:0 {0}(609,267)(585,267)(585,267)(562,267){1}
wire w174;    //: /sn:0 {0}(2213,425)(2152,425){1}
wire w20;    //: /sn:0 {0}(337,247)(326,247)(326,247)(316,247){1}
wire w23;    //: /sn:0 {0}(367,210)(396,210)(396,215)(460,215){1}
wire w242;    //: /sn:0 {0}(3017,495)(2934,495)(2934,495)(3052,495){1}
wire w108;    //: /sn:0 {0}(1098,318)(1103,318)(1103,318)(1110,318){1}
wire w225;    //: /sn:0 {0}(3207,482)(3219,482)(3219,480)(3237,480){1}
wire w82;    //: /sn:0 {0}(25,637)(2498,637)(2498,462){1}
//: {2}(2500,460)(2510,460)(2510,460)(2523,460){3}
//: {4}(2498,458)(2498,448)(2498,448)(2498,446)(2510,446)(2510,446)(2523,446){5}
wire w223;    //: /sn:0 {0}(2582,441)(2547,441)(2547,441)(2553,441){1}
wire w158;    //: /sn:0 {0}(1548,305)(1486,305){1}
wire w74;    //: /sn:0 {0}(25,567)(2035,567)(2035,427){1}
//: {2}(2037,425)(2047,425)(2047,425)(2060,425){3}
//: {4}(2035,423)(2035,413)(2035,413)(2035,399){5}
//: {6}(2037,397)(2060,397){7}
//: {8}(2035,395)(2035,388)(2035,388)(2035,375)(2035,375)(2035,355)(2060,355){9}
wire w91;    //: /sn:0 {0}(25,687)(2792,687)(2792,487){1}
//: {2}(2794,485)(2804,485)(2804,485)(2817,485){3}
//: {4}(2792,483)(2792,473)(2792,473)(2792,473){5}
//: {6}(2794,471)(2804,471)(2804,471)(2817,471){7}
//: {8}(2792,469)(2792,448)(2792,448)(2792,445){9}
//: {10}(2794,443)(2805,443)(2805,443)(2817,443){11}
//: {12}(2792,441)(2792,435)(2792,435)(2792,415)(2817,415){13}
wire w35;    //: /sn:0 {0}(609,253)(584,253)(584,253)(562,253){1}
wire w103;    //: /sn:0 {0}(987,277)(1051,277)(1051,294)(1112,294){1}
wire w8;    //: /sn:0 {0}(25,227)(179,227)(179,230){1}
//: {2}(181,228)(190,228)(190,228)(200,228){3}
//: {4}(179,226)(179,221)(179,221)(179,212){5}
//: {6}(181,214)(201,214){7}
//: {8}(179,216)(179,200)(201,200){9}
wire w192;    //: /sn:0 {0}(2339,435)(2291,435)(2291,435)(2307,435){1}
wire w163;    //: /sn:0 {0}(2122,420)(2087,420)(2087,420)(2090,420){1}
wire w101;    //: /sn:0 {0}(875,283)(883,283)(883,283)(894,283){1}
wire w238;    //: /sn:0 {0}(2938,429)(2889,429)(2889,429)(2908,429){1}
wire w202;    //: /sn:0 {0}(2339,407)(2291,407)(2291,407)(2307,407){1}
wire w71;    //: /sn:0 {0}(894,311)(888,311)(888,311)(875,311){1}
wire w144;    //: /sn:0 {0}(1392,338)(1368,338)(1368,338)(1345,338){1}
wire w22;    //: /sn:0 {0}(32,116)(32,157)(25,157){1}
wire w17;    //: /sn:0 {0}(269,242)(286,242){1}
wire w53;    //: /sn:0 {0}(25,407)(1060,407)(1060,338){1}
//: {2}(1062,336)(1067,336)(1067,336)(1068,336){3}
//: {4}(1060,334)(1060,325){5}
//: {6}(1062,323)(1065,323)(1065,323)(1068,323){7}
//: {8}(1060,321)(1060,288)(1070,288){9}
wire w84;    //: /sn:0 {0}(25,667)(2668,667)(2668,477){1}
//: {2}(2670,475)(2680,475)(2680,475)(2693,475){3}
//: {4}(2668,473)(2668,463)(2668,463)(2668,463){5}
//: {6}(2670,461)(2680,461)(2680,461)(2693,461){7}
//: {8}(2668,459)(2668,438)(2668,438)(2668,425)(2668,425)(2668,421){9}
//: {10}(2670,419)(2683,419)(2683,419)(2693,419){11}
//: {12}(2668,417)(2668,405)(2693,405){13}
wire w172;    //: /sn:0 {0}(1702,320)(1738,320)(1738,325)(1805,325){1}
wire w211;    //: /sn:0 {0}(2461,417)(2434,417)(2434,417)(2431,417){1}
wire w255;    //: /sn:0 {0}(3017,467)(3027,467)(3027,482)(2934,482)(2934,467)(3052,467){1}
wire w263;    //: /sn:0 {0}(3082,430)(3167,430)(3167,435)(3177,435){1}
wire w228;    //: /sn:0 {0}(2693,451)(2658,451)(2658,451)(2672,451){1}
wire w12;    //: /sn:0 {0}(147,179)(174,179)(174,190)(201,190){1}
wire w113;    //: /sn:0 {0}(1177,323)(1157,323)(1157,323)(1140,323){1}
wire w2;    //: /sn:0 {0}(78,172)(88,172)(88,174)(117,174){1}
wire w44;    //: /sn:0 {0}(705,291)(696,291)(696,291)(686,291){1}
wire w226;    //: /sn:0 {0}(2612,390)(2643,390)(2643,395)(2693,395){1}
wire w115;    //: /sn:0 {0}(1486,361)(1496,361)(1496,468)(2485,468)(2485,436)(2523,436){1}
wire w77;    //: /sn:0 {0}(25,617)(2376,617)(2376,452){1}
//: {2}(2378,450)(2388,450)(2388,450)(2401,450){3}
//: {4}(2376,448)(2376,438)(2376,438)(2376,424){5}
//: {6}(2378,422)(2401,422){7}
//: {8}(2376,420)(2376,413)(2376,413)(2376,410){9}
//: {10}(2378,408)(2389,408)(2389,408)(2401,408){11}
//: {12}(2376,406)(2376,400)(2376,400)(2376,394)(2391,394)(2391,394)(2401,394){13}
wire w83;    //: /sn:0 {0}(25,657)(2617,657)(2617,472){1}
//: {2}(2619,470)(2629,470)(2629,470)(2642,470){3}
//: {4}(2617,468)(2617,458)(2617,458)(2617,458){5}
//: {6}(2619,456)(2629,456)(2629,456)(2642,456){7}
//: {8}(2617,454)(2617,433)(2617,433)(2617,420)(2617,420)(2617,414)(2632,414)(2632,414)(2642,414){9}
wire w200;    //: /sn:0 {0}(2339,393)(2291,393)(2291,393)(2307,393){1}
wire w78;    //: /sn:0 {0}(779,245)(809,245)(809,248)(843,248){1}
wire w224;    //: /sn:0 {0}(2612,446)(2604,446)(2604,446)(2642,446){1}
wire w10;    //: /sn:0 {0}(318,219)(328,219)(328,219)(337,219){1}
wire w27;    //: /sn:0 {0}(230,223)(264,223)(264,238)(402,238){1}
wire w257;    //: /sn:0 {0}(3017,481)(2934,481)(2934,481)(3052,481){1}
wire w246;    //: /sn:0 {0}(2938,471)(2889,471)(2889,471)(2908,471){1}
wire w138;    //: /sn:0 {0}(1315,319)(1295,319)(1295,319)(1278,319){1}
wire w86;    //: /sn:0 {0}(25,647)(2557,647)(2557,467){1}
//: {2}(2559,465)(2569,465)(2569,465)(2582,465){3}
//: {4}(2557,463)(2557,453)(2557,453)(2557,453){5}
//: {6}(2559,451)(2569,451)(2569,451)(2582,451){7}
//: {8}(2557,449)(2557,428)(2557,428)(2557,415)(2557,415)(2557,395)(2582,395){9}
wire w188;    //: /sn:0 {0}(1964,354)(1998,354)(1998,364)(2122,364){1}
wire w52;    //: /sn:0 {0}(1046,313)(1056,313)(1056,313)(1068,313){1}
wire w95;    //: /sn:0 {0}(25,707)(2913,707)(2913,497){1}
//: {2}(2915,495)(2925,495)(2925,495)(2938,495){3}
//: {4}(2913,493)(2913,483)(2913,483)(2913,483){5}
//: {6}(2915,481)(2925,481)(2925,481)(2938,481){7}
//: {8}(2913,479)(2913,458)(2913,458)(2913,455){9}
//: {10}(2915,453)(2926,453)(2926,453)(2938,453){11}
//: {12}(2913,451)(2913,445)(2913,445)(2913,441){13}
//: {14}(2915,439)(2928,439)(2928,439)(2938,439){15}
//: {16}(2913,437)(2913,425)(2938,425){17}
wire w231;    //: /sn:0 {0}(2817,433)(2785,433)(2785,433)(2784,433){1}
wire w29;    //: /sn:0 {0}(25,187)(38,187){1}
//: {2}(40,185)(40,177)(48,177){3}
//: {4}(40,189)(40,193)(55,193){5}
wire w80;    //: /sn:0 {0}(25,597)(2252,597)(2252,442){1}
//: {2}(2254,440)(2264,440)(2264,440)(2277,440){3}
//: {4}(2252,438)(2252,428)(2252,428)(2252,414){5}
//: {6}(2254,412)(2277,412){7}
//: {8}(2252,410)(2252,403)(2252,403)(2252,398)(2265,398)(2265,398)(2277,398){9}
wire w155;    //: /sn:0 {0}(2020,387)(2021,387)(2021,387)(2060,387){1}
wire w178;    //: /sn:0 {0}(1934,335)(1913,335)(1913,330)(1835,330){1}
wire w142;    //: /sn:0 {0}(1278,346)(1285,346)(1285,346)(1317,346){1}
wire w147;    //: /sn:0 {0}(1317,290)(1230,290)(1230,290)(1207,290){1}
wire w42;    //: /sn:0 {0}(461,253)(454,253)(454,253)(447,253){1}
//: {2}(445,251)(445,225)(460,225){3}
//: {4}(445,255)(445,271)(445,271)(445,269){5}
//: {6}(447,267)(454,267)(454,267)(461,267){7}
//: {8}(443,267)(433,267)(433,287)(25,287){9}
wire w50;    //: /sn:0 {0}(845,288)(834,288){1}
//: {2}(832,286)(832,258)(843,258){3}
//: {4}(832,290)(832,314){5}
//: {6}(834,316)(840,316)(840,316)(845,316){7}
//: {8}(832,318)(832,367)(25,367){9}
wire w6;    //: /sn:0 {0}(25,197)(85,197)(85,201)(116,201){1}
wire w247;    //: /sn:0 {0}(2968,448)(3099,448)(3099,470)(3237,470){1}
wire w7;    //: /sn:0 {0}(25,217)(130,217)(130,223)(140,223){1}
//: {2}(144,223)(158,223){3}
//: {4}(142,221)(142,209)(158,209){5}
wire w93;    //: /sn:0 {0}(25,677)(2729,677)(2729,482){1}
//: {2}(2731,480)(2741,480)(2741,480)(2754,480){3}
//: {4}(2729,478)(2729,468)(2729,468)(2729,468){5}
//: {6}(2731,466)(2741,466)(2741,466)(2754,466){7}
//: {8}(2729,464)(2729,443)(2729,443)(2729,438)(2742,438)(2742,438)(2754,438){9}
wire w175;    //: /sn:0 {0}(1934,363)(1883,363)(1883,363)(1902,363){1}
wire w112;    //: /sn:0 {0}(3207,454)(3219,454)(3219,460)(3237,460){1}
wire w46;    //: /sn:0 {0}(686,235)(705,235)(705,240)(749,240){1}
wire w60;    //: /sn:0 {0}(25,477)(1480,477)(1480,375)(1548,375){1}
wire w99;    //: /sn:0 {0}(924,272)(937,272)(937,272)(957,272){1}
wire w61;    //: /sn:0 {0}(25,277)(385,277)(385,264){1}
//: {2}(387,262)(397,262)(397,262)(402,262){3}
//: {4}(385,260)(385,248)(402,248){5}
wire w153;    //: /sn:0 {0}(1702,390)(1695,390)(1695,390)(1730,390){1}
wire w135;    //: /sn:0 {0}(1392,324)(1367,324)(1367,324)(1345,324){1}
wire w15;    //: /sn:0 {0}(188,204)(191,204)(191,204)(201,204){1}
wire w216;    //: /sn:0 {0}(2693,465)(2658,465)(2658,465)(2672,465){1}
wire w207;    //: /sn:0 {0}(2642,460)(2604,460)(2604,460)(2612,460){1}
wire w239;    //: /sn:0 {0}(2987,490)(2968,490){1}
wire w109;    //: /sn:0 {0}(1111,331)(1100,331)(1100,331)(1098,331){1}
wire w51;    //: /sn:0 {0}(894,321)(888,321)(888,321)(880,321){1}
//: {2}(878,319)(878,295){3}
//: {4}(880,293)(888,293)(888,293)(894,293){5}
//: {6}(878,291)(878,277)(894,277){7}
//: {8}(878,323)(878,377)(25,377){9}
wire w69;    //: /sn:0 {0}(25,447)(1292,447)(1292,358){1}
//: {2}(1294,356)(1304,356)(1304,356)(1317,356){3}
//: {4}(1292,354)(1292,349)(1292,349)(1292,345){5}
//: {6}(1294,343)(1304,343)(1304,343)(1315,343){7}
//: {8}(1292,341)(1292,331){9}
//: {10}(1294,329)(1303,329)(1303,329)(1315,329){11}
//: {12}(1292,327)(1292,300)(1317,300){13}
wire w213;    //: /sn:0 {0}(2491,408)(2520,408)(2520,416)(2608,416)(2608,428)(2754,428){1}
wire w229;    //: /sn:0 {0}(2878,480)(2826,480)(2826,480)(2847,480){1}
wire w114;    //: /sn:0 {0}(2369,398)(2364,398)(2364,398)(2401,398){1}
wire w97;    //: /sn:0 {0}(25,717)(2975,717)(2975,502){1}
//: {2}(2977,500)(2987,500)(2987,500)(2987,500){3}
//: {4}(2975,498)(2975,488)(2975,488)(2975,488){5}
//: {6}(2977,486)(2987,486)(2987,486)(2987,486){7}
//: {8}(2975,484)(2975,472)(2987,472){9}
wire w245;    //: /sn:0 {0}(2908,443)(2889,443)(2889,443)(2938,443){1}
wire w64;    //: /sn:0 {0}(656,296)(656,296)(656,296)(646,296){1}
//: {2}(644,294)(644,240)(656,240){3}
//: {4}(644,298)(644,327)(25,327){5}
wire w261;    //: /sn:0 {0}(3082,486)(3075,486)(3075,486)(3114,486){1}
wire w177;    //: /sn:0 {0}(2213,369)(2152,369){1}
wire w66;    //: /sn:0 {0}(1835,400)(1823,400)(1823,400)(1872,400){1}
wire w37;    //: /sn:0 {0}(609,239)(582,239)(582,239)(562,239){1}
wire w159;    //: /sn:0 {0}(2060,415)(2023,415)(2023,415)(2020,415){1}
wire w63;    //: /sn:0 {0}(1612,390)(1599,390)(1599,390)(1589,390){1}
//: {2}(1587,388)(1587,378)(1587,378)(1587,353)(1587,353)(1587,340)(1587,340)(1587,334)(1602,334)(1602,334)(1612,334){3}
//: {4}(1587,392)(1587,497)(25,497){5}
wire w259;    //: /sn:0 {0}(3082,472)(3075,472)(3075,472)(3114,472){1}
wire w234;    //: /sn:0 {0}(2723,400)(2793,400)(2793,405)(2817,405){1}
wire w34;    //: /sn:0 {0}(639,230)(640,230)(640,230)(656,230){1}
wire w236;    //: /sn:0 {0}(2878,438)(2826,438)(2826,438)(2847,438){1}
wire w21;    //: /sn:0 {0}(432,243)(455,243)(455,243)(461,243){1}
wire w76;    //: /sn:0 {0}(25,577)(2097,577)(2097,432){1}
//: {2}(2099,430)(2109,430)(2109,430)(2122,430){3}
//: {4}(2097,428)(2097,418)(2097,418)(2097,404){5}
//: {6}(2099,402)(2122,402){7}
//: {8}(2097,400)(2097,393)(2097,393)(2097,380)(2097,380)(2097,374)(2112,374)(2112,374)(2122,374){9}
wire w157;    //: /sn:0 {0}(1612,380)(1576,380)(1576,380)(1578,380){1}
wire w102;    //: /sn:0 {0}(924,316)(937,316)(937,316)(957,316){1}
wire w43;    //: /sn:0 {0}(367,224)(424,224)(424,234)(532,234){1}
wire w87;    //: /sn:0 {0}(796,301)(779,301){1}
wire w199;    //: /sn:0 {0}(2339,365)(2317,365)(2317,360)(2243,360){1}
wire w170;    //: /sn:0 {0}(1964,410)(1938,410)(1938,410)(1990,410){1}
wire w100;    //: /sn:0 {0}(25,727)(3027,727)(3027,507){1}
//: {2}(3029,505)(3039,505)(3039,505)(3052,505){3}
//: {4}(3027,503)(3027,493)(3027,493)(3027,493){5}
//: {6}(3029,491)(3039,491)(3039,491)(3052,491){7}
//: {8}(3027,489)(3027,479){9}
//: {10}(3029,477)(3052,477){11}
//: {12}(3027,475)(3027,468)(3027,468)(3027,455)(3027,455)(3027,435)(3052,435){13}
wire w31;    //: /sn:0 {0}(749,254)(738,254)(738,254)(736,254){1}
wire w249;    //: /sn:0 {0}(3082,500)(3075,500)(3075,500)(3114,500){1}
wire w58;    //: /sn:0 {0}(1392,361)(1380,361)(1380,361)(1369,361){1}
//: {2}(1367,359)(1367,355)(1367,355)(1367,350){3}
//: {4}(1369,348)(1380,348)(1380,348)(1392,348){5}
//: {6}(1367,346)(1367,341)(1367,341)(1367,336){7}
//: {8}(1369,334)(1380,334)(1380,334)(1392,334){9}
//: {10}(1367,332)(1367,321)(1392,321){11}
//: {12}(1367,363)(1367,457)(25,457){13}
wire w169;    //: /sn:0 {0}(1902,405)(1883,405)(1883,405)(1934,405){1}
wire w130;    //: /sn:0 {0}(987,321)(997,321)(997,321)(1016,321){1}
wire w28;    //: /sn:0 {0}(25,177)(37,177)(37,183)(55,183){1}
wire w251;    //: /sn:0 {0}(2987,476)(2971,476)(2971,476)(2968,476){1}
wire w161;    //: /sn:0 {0}(1702,334)(1739,334)(1739,344)(1872,344){1}
wire w132;    //: /sn:0 {0}(367,252)(397,252)(397,252)(402,252){1}
wire w1;    //: /sn:0 {0}(1068,326)(1058,326)(1058,326)(1046,326){1}
wire w241;    //: /sn:0 {0}(2878,466)(2826,466)(2826,466)(2847,466){1}
wire w140;    //: /sn:0 {0}(1278,333)(1296,333)(1296,333)(1315,333){1}
wire w235;    //: /sn:0 {0}(3207,496)(3216,496)(3216,490)(3237,490){1}
wire w253;    //: /sn:0 {0}(3052,425)(3028,425)(3028,420)(2968,420){1}
wire w205;    //: /sn:0 {0}(2461,389)(2434,389)(2434,389)(2431,389){1}
wire w154;    //: /sn:0 {0}(1642,329)(1649,329)(1649,329)(1672,329){1}
wire w25;    //: /sn:0 {0}(25,167)(48,167){1}
wire w227;    //: /sn:0 {0}(2784,475)(2776,475)(2776,475)(2817,475){1}
wire w116;    //: /sn:0 {0}(1177,299)(1166,299)(1166,299)(1142,299){1}
wire w98;    //: /sn:0 {0}(845,306)(836,306)(836,306)(826,306){1}
wire w210;    //: /sn:0 {0}(2461,375)(2453,375)(2453,370)(2369,370){1}
wire w65;    //: /sn:0 {0}(25,507)(1647,507)(1647,397){1}
//: {2}(1649,395)(1659,395)(1659,395)(1672,395){3}
//: {4}(1647,393)(1647,358)(1647,358)(1647,341){5}
//: {6}(1649,339)(1672,339){7}
//: {8}(1647,337)(1647,325)(1672,325){9}
wire w243;    //: /sn:0 {0}(2938,415)(2912,415)(2912,410)(2847,410){1}
wire w212;    //: /sn:0 {0}(2582,455)(2547,455)(2547,455)(2553,455){1}
wire w18;    //: /sn:0 {0}(25,237)(210,237)(210,237)(239,237){1}
wire w40;    //: /sn:0 {0}(25,307)(578,307)(578,277)(588,277){1}
//: {2}(592,277)(601,277)(601,277)(609,277){3}
//: {4}(590,279)(590,280)(590,280)(590,265){5}
//: {6}(592,263)(593,263)(593,263)(609,263){7}
//: {8}(590,261)(590,253)(590,253)(590,251){9}
//: {10}(592,249)(599,249)(599,249)(609,249){11}
//: {12}(590,247)(590,235)(609,235){13}
wire w92;    //: /sn:0 {0}(845,278)(834,278)(834,278)(824,278){1}
wire w164;    //: /sn:0 {0}(1486,334)(1507,334)(1507,348)(1730,348){1}
wire w68;    //: /sn:0 {0}(1805,405)(1792,405)(1792,405)(1782,405){1}
//: {2}(1780,403)(1780,393)(1780,393)(1780,368)(1780,368)(1780,365){3}
//: {4}(1782,363)(1793,363)(1793,363)(1805,363){5}
//: {6}(1780,361)(1780,355)(1780,355)(1780,335)(1805,335){7}
//: {8}(1780,407)(1780,527)(25,527){9}
wire w162;    //: /sn:0 {0}(1760,395)(1759,395)(1759,395)(1805,395){1}
wire w30;    //: /sn:0 {0}(432,257)(436,257)(436,257)(461,257){1}
wire w198;    //: /sn:0 {0}(3144,477)(3142,477)(3142,477)(3177,477){1}
wire w222;    //: /sn:0 {0}(2723,414)(2734,414)(2734,424)(2878,424){1}
wire w149;    //: /sn:0 {0}(1964,340)(2037,340)(2037,345)(2060,345){1}
wire w146;    //: /sn:0 {0}(1392,351)(1357,351)(1357,351)(1347,351){1}
wire w59;    //: /sn:0 {0}(25,467)(1431,467)(1431,368){1}
//: {2}(1433,366)(1443,366)(1443,366)(1456,366){3}
//: {4}(1431,364)(1431,360)(1431,360)(1431,355){5}
//: {6}(1433,353)(1444,353)(1444,353)(1456,353){7}
//: {8}(1431,351)(1431,346)(1431,346)(1431,341){9}
//: {10}(1433,339)(1444,339)(1444,339)(1456,339){11}
//: {12}(1431,337)(1431,333)(1431,333)(1431,328){13}
//: {14}(1433,326)(1444,326)(1444,326)(1456,326){15}
//: {16}(1431,324)(1431,310)(1456,310){17}
wire w62;    //: /sn:0 {0}(25,487)(1523,487)(1523,387){1}
//: {2}(1525,385)(1535,385)(1535,385)(1548,385){3}
//: {4}(1523,383)(1523,373)(1523,373)(1523,348)(1523,348)(1523,335)(1523,335)(1523,315)(1548,315){5}
wire w85;    //: /sn:0 {0}(749,296)(736,296)(736,296)(735,296){1}
wire w248;    //: /sn:0 {0}(3207,440)(3217,440)(3217,450)(3237,450){1}
wire w197;    //: /sn:0 {0}(2401,440)(2364,440)(2364,440)(2369,440){1}
wire w137;    //: /sn:0 {0}(1207,341)(1244,341)(1244,341)(1248,341){1}
wire w11;    //: /sn:0 {0}(337,229)(331,229)(331,229)(325,229){1}
//: {2}(323,227)(323,215)(337,215){3}
//: {4}(323,231)(323,243)(323,243)(323,255){5}
//: {6}(325,257)(330,257)(330,257)(337,257){7}
//: {8}(323,259)(323,267)(25,267){9}
wire w173;    //: /sn:0 {0}(1934,349)(1883,349)(1883,349)(1902,349){1}
wire w139;    //: /sn:0 {0}(25,517)(1705,517)(1705,402){1}
//: {2}(1707,400)(1717,400)(1717,400)(1730,400){3}
//: {4}(1705,398)(1705,388)(1705,388)(1705,363)(1705,363)(1705,358)(1718,358)(1718,358)(1730,358){5}
wire w57;    //: /sn:0 {0}(1612,324)(1553,324)(1553,321)(1486,321){1}
wire w136;    //: /sn:0 {0}(1456,329)(1439,329)(1439,329)(1422,329){1}
wire w49;    //: /sn:0 {0}(794,273)(704,273)(704,267)(653,267)(653,258)(639,258){1}
wire w189;    //: /sn:0 {0}(2213,397)(2152,397){1}
wire w150;    //: /sn:0 {0}(1456,343)(1439,343)(1439,343)(1422,343){1}
wire w110;    //: /sn:0 {0}(1141,336)(1169,336)(1169,336)(1177,336){1}
wire w70;    //: /sn:0 {0}(1872,410)(1859,410)(1859,410)(1849,410){1}
//: {2}(1847,408)(1847,398)(1847,398)(1847,373)(1847,373)(1847,370){3}
//: {4}(1849,368)(1860,368)(1860,368)(1872,368){5}
//: {6}(1847,366)(1847,360)(1847,360)(1847,354)(1862,354)(1862,354)(1872,354){7}
//: {8}(1847,412)(1847,537)(25,537){9}
wire w193;    //: /sn:0 {0}(1934,415)(1921,415)(1921,415)(1911,415){1}
//: {2}(1909,413)(1909,403)(1909,403)(1909,378)(1909,378)(1909,375){3}
//: {4}(1911,373)(1922,373)(1922,373)(1934,373){5}
//: {6}(1909,371)(1909,365)(1910,365)(1910,361){7}
//: {8}(1912,359)(1934,359){9}
//: {10}(1910,357)(1910,345)(1934,345){11}
//: {12}(1909,417)(1909,547)(25,547){13}
wire w148;    //: /sn:0 {0}(1422,356)(1456,356){1}
wire w105;    //: /sn:0 {0}(1964,368)(2010,368)(2010,376)(2042,376)(2042,382)(2136,382)(2136,388)(2277,388){1}
wire w206;    //: /sn:0 {0}(2401,412)(2364,412)(2364,412)(2369,412){1}
wire w13;    //: /sn:0 {0}(146,196)(152,196)(152,213)(158,213){1}
wire w88;    //: /sn:0 {0}(779,259)(825,259)(825,267)(894,267){1}
wire w94;    //: /sn:0 {0}(957,326)(947,326)(947,326)(944,326){1}
//: {2}(942,324)(942,317)(942,317)(942,300){3}
//: {4}(944,298)(951,298)(951,298)(957,298){5}
//: {6}(942,296)(942,287)(942,287)(942,284){7}
//: {8}(944,282)(951,282)(951,282)(957,282){9}
//: {10}(942,280)(942,268)(957,268){11}
//: {12}(942,328)(942,387)(25,387){13}
wire w72;    //: /sn:0 {0}(25,587)(2188,587)(2188,437){1}
//: {2}(2190,435)(2200,435)(2200,435)(2213,435){3}
//: {4}(2188,433)(2188,423)(2188,423)(2188,409){5}
//: {6}(2190,407)(2213,407){7}
//: {8}(2188,405)(2188,398)(2188,398)(2188,385)(2188,385)(2188,381){9}
//: {10}(2190,379)(2203,379)(2203,379)(2213,379){11}
//: {12}(2188,377)(2188,365)(2213,365){13}
wire w208;    //: /sn:0 {0}(2431,403)(2434,403)(2434,403)(2461,403){1}
wire w5;    //: /sn:0 {0}(271,200)(280,200)(280,205)(337,205){1}
wire w48;    //: /sn:0 {0}(794,283)(785,283)(785,309){1}
//: {2}(787,311)(796,311){3}
//: {4}(785,313)(785,357)(25,357){5}
wire w33;    //: /sn:0 {0}(532,248)(504,248)(504,248)(491,248){1}
wire w191;    //: /sn:0 {0}(3207,510)(3218,510)(3218,500)(3237,500){1}
wire w47;    //: /sn:0 {0}(749,264)(745,264)(745,264)(742,264){1}
//: {2}(740,262)(740,250)(749,250){3}
//: {4}(740,266)(740,304){5}
//: {6}(742,306)(744,306)(744,306)(749,306){7}
//: {8}(740,308)(740,347)(25,347){9}
wire w143;    //: /sn:0 {0}(1486,348)(1489,348)(1489,358)(1702,358)(1702,382)(1990,382){1}
wire w107;    //: /sn:0 {0}(1100,283)(1167,283)(1167,285)(1177,285){1}
wire w219;    //: /sn:0 {0}(2491,380)(2558,380)(2558,385)(2582,385){1}
wire w9;    //: /sn:0 {0}(25,207)(101,207)(101,193){1}
//: {2}(103,191)(116,191){3}
//: {4}(101,189)(101,184)(117,184){5}
wire w79;    //: /sn:0 {0}(25,607)(2314,607)(2314,447){1}
//: {2}(2316,445)(2326,445)(2326,445)(2339,445){3}
//: {4}(2314,443)(2314,433)(2314,433)(2314,419){5}
//: {6}(2316,417)(2339,417){7}
//: {8}(2314,415)(2314,408)(2314,408)(2314,405){9}
//: {10}(2316,403)(2327,403)(2327,403)(2339,403){11}
//: {12}(2314,401)(2314,395)(2314,395)(2314,375)(2339,375){13}
wire w232;    //: /sn:0 {0}(2723,456)(2710,456)(2710,456)(2754,456){1}
wire w201;    //: /sn:0 {0}(2461,445)(2434,445)(2434,445)(2431,445){1}
wire w55;    //: /sn:0 {0}(25,417)(1098,417)(1098,343){1}
//: {2}(1100,341)(1105,341)(1105,341)(1111,341){3}
//: {4}(1098,339)(1098,335)(1098,335)(1098,330){5}
//: {6}(1100,328)(1104,328)(1104,328)(1110,328){7}
//: {8}(1098,326)(1098,304)(1112,304){9}
wire w39;    //: /sn:0 {0}(957,288)(940,288)(940,288)(924,288){1}
//: enddecls

  OrMos g8 (.A(w5), .B(w11), .Z(w23));   //: @(353, 210) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g165 (w68) @(1780, 363) /w:[ 4 6 -1 3 ]
  //: joint g55 (w64) @(644, 296) /w:[ 1 2 -1 4 ]
  //: joint g13 (w9) @(101, 191) /w:[ 2 4 -1 1 ]
  //: joint g37 (w42) @(445, 253) /w:[ 1 2 -1 4 ]
  //: joint g111 (w133) @(1223, 338) /w:[ 6 8 -1 5 ]
  //: joint g176 (w74) @(2035, 397) /w:[ 6 8 -1 5 ]
  OrMos g218 (.A(w204), .B(w82), .Z(w212));   //: @(2539, 455) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g1 (.A(w2), .B(w9), .Z(w12));   //: @(133, 179) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g277 (.A(w249), .B(w96), .Z(w166));   //: @(3130, 505) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g11 (.A(w4), .B(w7), .Z(w15));   //: @(174, 204) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g130 (.A(w151), .B(w58), .Z(w152));   //: @(1408, 316) /symbol:3101448544 /sn:0 /w:[ 1 11 1 ]
  //: joint g266 (w95) @(2913, 481) /w:[ 6 8 -1 5 ]
  OrMos g50 (.A(w25), .B(w29), .Z(w2));   //: @(64, 172) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g254 (.A(w234), .B(w91), .Z(w243));   //: @(2833, 410) /symbol:3101448544 /sn:0 /w:[ 1 13 1 ]
  OrMos g306 (.A(w20), .B(w11), .Z(w132));   //: @(353, 252) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g113 (.A(w134), .B(w133), .Z(w138));   //: @(1264, 319) /symbol:3101448544 /sn:0 /w:[ 0 9 1 ]
  //: joint g19 (w8) @(179, 214) /w:[ 6 5 -1 8 ]
  OrMos g132 (.A(w136), .B(w59), .Z(w164));   //: @(1472, 334) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  OrMos g197 (.A(w195), .B(w80), .Z(w202));   //: @(2293, 407) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g223 (.A(w212), .B(w86), .Z(w207));   //: @(2598, 460) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g150 (.A(w158), .B(w62), .Z(w168));   //: @(1564, 310) /symbol:3101448544 /sn:0 /w:[ 0 5 0 ]
  OrMos g146 (.A(w57), .B(w63), .Z(w154));   //: @(1628, 329) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  //: joint g115 (w133) @(1223, 351) /w:[ 2 4 -1 1 ]
  OrMos g38 (.A(w43), .B(w156), .Z(w37));   //: @(548, 239) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  //: joint g307 (w11) @(323, 257) /w:[ 6 5 -1 8 ]
  OrMos g75 (.A(w104), .B(w94), .Z(w89));   //: @(973, 263) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  OrMos g20 (.A(w12), .B(w8), .Z(w16));   //: @(217, 195) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  //: joint g135 (w59) @(1431, 366) /w:[ 2 4 -1 1 ]
  //: joint g160 (w193) @(1909, 415) /w:[ 1 2 -1 12 ]
  OrMos g169 (.A(w170), .B(w75), .Z(w159));   //: @(2006, 415) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  //: joint g227 (w84) @(2668, 475) /w:[ 2 4 -1 1 ]
  //: joint g31 (w94) @(942, 326) /w:[ 1 2 -1 12 ]
  //: joint g124 (w69) @(1292, 329) /w:[ 10 12 -1 9 ]
  //: joint g230 (w86) @(2557, 451) /w:[ 6 8 -1 5 ]
  OrMos g68 (.A(w98), .B(w50), .Z(w71));   //: @(861, 311) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  //: joint g39 (w42) @(445, 267) /w:[ 6 -1 8 5 ]
  //: joint g284 (w41) @(3152, 515) /w:[ 2 4 -1 1 ]
  //: joint g195 (w79) @(2314, 445) /w:[ 2 4 -1 1 ]
  //: joint g52 (w40) @(590, 277) /w:[ 2 -1 1 4 ]
  OrMos g179 (.A(w163), .B(w76), .Z(w174));   //: @(2138, 425) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g205 (.A(w182), .B(w77), .Z(w205));   //: @(2417, 389) /symbol:3101448544 /sn:0 /w:[ 1 13 1 ]
  OrMos g231 (.A(w216), .B(w84), .Z(w220));   //: @(2709, 470) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  OrMos g201 (.A(w200), .B(w79), .Z(w114));   //: @(2355, 398) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  //: joint g221 (w81) @(2436, 413) /w:[ 10 12 -1 9 ]
  OrMos g14 (.A(w23), .B(w42), .Z(w45));   //: @(476, 220) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g44 (.A(w45), .B(w40), .Z(w34));   //: @(625, 230) /symbol:3101448544 /sn:0 /w:[ 1 13 0 ]
  OrMos g47 (.A(w35), .B(w40), .Z(w49));   //: @(625, 258) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  OrMos g84 (.A(w1), .B(w53), .Z(w109));   //: @(1084, 331) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  //: joint g247 (w93) @(2729, 466) /w:[ 6 8 -1 5 ]
  OrMos g236 (.A(w218), .B(w84), .Z(w222));   //: @(2709, 414) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  //: joint g23 (w61) @(385, 262) /w:[ 2 4 -1 1 ]
  OrMos g116 (.A(w137), .B(w133), .Z(w142));   //: @(1264, 346) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g93 (w55) @(1098, 341) /w:[ 2 4 -1 1 ]
  OrMos g40 (.A(w33), .B(w156), .Z(w35));   //: @(548, 253) /symbol:3101448544 /sn:0 /w:[ 0 5 1 ]
  //: joint g54 (w29) @(40, 187) /w:[ -1 2 1 4 ]
  OrMos g249 (.A(w231), .B(w91), .Z(w236));   //: @(2833, 438) /symbol:3101448544 /sn:0 /w:[ 0 11 1 ]
  OrMos g26 (.A(w15), .B(w8), .Z(w0));   //: @(217, 209) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  //: comment g0 @(689,-183) /sn:0
  //: /line:"dec| bin |  my"
  //: /line:""
  //: /line:"00 | 000000 21 | 010101 42 | 101010 63 |  111111"
  //: /line:"01 | 000001 22 | 010110 43 | 101011 "
  //: /line:"02 | 000010 23 | 010111 44 | 101100"
  //: /line:"03 | 000011 24 | 011000 45 | 101101"
  //: /line:"04 | 000100 25 | 011001 46 | 101110"
  //: /line:"05 | 000101 26 | 011010 47 | 101111"
  //: /line:"06 | 000110 27 | 011011 48 | 110000"
  //: /line:"07 | 000111 28 | 011100 49 | 110001"
  //: /line:"08 | 001000 29 | 011101 50 | 110010"
  //: /line:"09 | 001001 30 | 011110 51 | 110011"
  //: /line:"10 | 001010 31 | 011111 52 | 110100"
  //: /line:"11 | 001011 32 | 100000 53 | 110101"
  //: /line:"12 | 001100 33 | 100001 54 | 110110"
  //: /line:"13 | 001101 34 | 100010 55 | 110111"
  //: /line:"14 | 001110 35 | 100011 56 | 111000"
  //: /line:"15 | 001111 36 | 100100 57 | 111001"
  //: /line:"16 | 010000 37 | 100101 58 | 111010"
  //: /line:"17 | 010001 38 | 100110 59 | 111011"
  //: /line:"18 | 010010 39 | 100111 60 | 111100"
  //: /line:"19 | 010011 40 | 101000 61 | 111101"
  //: /line:"20 | 010100 41 | 101001 62 | 111110"
  //: /line:""
  //: /end
  //: joint g46 (w40) @(590, 249) /w:[ 10 12 -1 9 ]
  OrMos g167 (.A(w173), .B(w193), .Z(w188));   //: @(1950, 354) /symbol:3101448544 /sn:0 /w:[ 0 9 0 ]
  OrMos g278 (.A(w255), .B(w100), .Z(w259));   //: @(3068, 472) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  OrMos g228 (.A(w209), .B(w83), .Z(w218));   //: @(2658, 409) /symbol:3101448544 /sn:0 /w:[ 0 9 1 ]
  //: joint g136 (w59) @(1431, 326) /w:[ 14 16 -1 13 ]
  //: joint g224 (w83) @(2617, 470) /w:[ 2 4 -1 1 ]
  //: joint g233 (w93) @(2729, 480) /w:[ 2 4 -1 1 ]
  //: joint g173 (w193) @(1910, 359) /w:[ 8 10 -1 7 ]
  OrMos g190 (.A(w189), .B(w72), .Z(w195));   //: @(2229, 402) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g61 (.A(w92), .B(w50), .Z(w101));   //: @(861, 283) /symbol:3101448544 /sn:0 /w:[ 0 0 0 ]
  OrMos g34 (.A(w19), .B(w64), .Z(w44));   //: @(672, 291) /symbol:3101448544 /sn:0 /w:[ 0 0 1 ]
  OrMos g3 (.A(w28), .B(w29), .Z(w4));   //: @(71, 188) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  //: joint g86 (w53) @(1060, 323) /w:[ 6 8 -1 5 ]
  OrMos g220 (.A(w210), .B(w81), .Z(w219));   //: @(2477, 380) /symbol:3101448544 /sn:0 /w:[ 0 17 0 ]
  //: joint g267 (w95) @(2913, 439) /w:[ 14 16 -1 13 ]
  OrMos g261 (.A(w238), .B(w95), .Z(w244));   //: @(2954, 434) /symbol:3101448544 /sn:0 /w:[ 0 15 0 ]
  //: joint g250 (w95) @(2913, 495) /w:[ 2 4 -1 1 ]
  OrMos g110 (.A(w130), .B(w54), .Z(w1));   //: @(1032, 326) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  OrMos g65 (.A(w87), .B(w48), .Z(w98));   //: @(812, 306) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  //: joint g59 (w67) @(693, 301) /w:[ 2 4 -1 1 ]
  OrMos g147 (.A(w160), .B(w65), .Z(w153));   //: @(1688, 390) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  OrMos g156 (.A(w168), .B(w65), .Z(w172));   //: @(1688, 320) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  OrMos g153 (.A(w162), .B(w68), .Z(w66));   //: @(1821, 400) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: joint g98 (w56) @(1153, 346) /w:[ 1 2 -1 12 ]
  //: joint g16 (w7) @(142, 223) /w:[ 2 4 1 -1 ]
  //: joint g96 (w56) @(1153, 309) /w:[ 8 10 -1 7 ]
  OrMos g122 (.A(w135), .B(w58), .Z(w136));   //: @(1408, 329) /symbol:3101448544 /sn:0 /w:[ 0 9 1 ]
  //: joint g183 (w72) @(2188, 435) /w:[ 2 4 -1 1 ]
  //: joint g280 (w100) @(3027, 491) /w:[ 6 8 -1 5 ]
  OrMos g87 (.A(w108), .B(w55), .Z(w113));   //: @(1126, 323) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  //: joint g78 (w53) @(1060, 336) /w:[ 2 4 -1 1 ]
  //: joint g129 (w58) @(1367, 334) /w:[ 8 10 -1 7 ]
  //: joint g171 (w74) @(2035, 425) /w:[ 2 4 -1 1 ]
  OrMos g258 (.A(w241), .B(w90), .Z(w246));   //: @(2894, 471) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  //: joint g69 (w50) @(832, 316) /w:[ 6 5 -1 8 ]
  //: joint g143 (w63) @(1587, 390) /w:[ 1 2 -1 4 ]
  OrMos g244 (.A(w213), .B(w93), .Z(w231));   //: @(2770, 433) /symbol:3101448544 /sn:0 /w:[ 1 9 1 ]
  //: joint g245 (w90) @(2853, 490) /w:[ 2 4 -1 1 ]
  OrMos g119 (.A(w140), .B(w69), .Z(w144));   //: @(1331, 338) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g15 (.A(w18), .B(w3), .Z(w17));   //: @(255, 242) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g162 (.A(w171), .B(w70), .Z(w175));   //: @(1888, 363) /symbol:3101448544 /sn:0 /w:[ 0 5 1 ]
  //: joint g67 (w50) @(832, 288) /w:[ 1 2 -1 4 ]
  //: joint g131 (w58) @(1367, 348) /w:[ 4 6 -1 3 ]
  //: joint g127 (w59) @(1431, 353) /w:[ 6 8 -1 5 ]
  OrMos g293 (.A(w176), .B(w41), .Z(w235));   //: @(3193, 496) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  //: joint g43 (w156) @(513, 272) /w:[ 1 2 -1 8 ]
  //: joint g62 (w47) @(740, 264) /w:[ 1 2 -1 4 ]
  OrMos g63 (.A(w85), .B(w47), .Z(w87));   //: @(765, 301) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  //: joint g138 (w59) @(1431, 339) /w:[ 10 12 -1 9 ]
  OrMos g188 (.A(w177), .B(w72), .Z(w182));   //: @(2229, 374) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  OrMos g257 (.A(w233), .B(w95), .Z(w239));   //: @(2954, 490) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  //: joint g109 (w54) @(998, 331) /w:[ 2 4 -1 1 ]
  //: joint g175 (w193) @(1909, 373) /w:[ 4 6 -1 3 ]
  OrMos g234 (.A(w224), .B(w83), .Z(w228));   //: @(2658, 451) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g285 (.A(w259), .B(w96), .Z(w198));   //: @(3130, 477) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  OrMos g264 (.A(w239), .B(w97), .Z(w242));   //: @(3003, 495) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  OrMos g56 (.A(w34), .B(w64), .Z(w46));   //: @(672, 235) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: IN g5 (pos) @(-27,452) /sn:0 /w:[ 0 ]
  OrMos g133 (.A(w150), .B(w59), .Z(w143));   //: @(1472, 348) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  //: joint g95 (w56) @(1153, 333) /w:[ 4 6 -1 3 ]
  OrMos g24 (.A(w27), .B(w61), .Z(w21));   //: @(418, 243) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g85 (.A(w109), .B(w55), .Z(w110));   //: @(1127, 336) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  OrMos g92 (.A(w116), .B(w56), .Z(w151));   //: @(1193, 304) /symbol:3101448544 /sn:0 /w:[ 0 9 0 ]
  //: joint g210 (w81) @(2436, 455) /w:[ 2 4 -1 1 ]
  OrMos g60 (.A(w49), .B(w48), .Z(w92));   //: @(810, 278) /symbol:3101448544 /sn:0 /w:[ 0 0 1 ]
  //: joint g214 (w77) @(2376, 408) /w:[ 10 12 -1 9 ]
  OrMos g185 (.A(w179), .B(w76), .Z(w189));   //: @(2138, 397) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  //: joint g170 (w70) @(1847, 368) /w:[ 4 6 -1 3 ]
  OrMos g126 (.A(w146), .B(w58), .Z(w148));   //: @(1408, 356) /symbol:3101448544 /sn:0 /w:[ 0 0 0 ]
  OrMos g35 (.A(w73), .B(w67), .Z(w31));   //: @(722, 254) /symbol:3101448544 /sn:0 /w:[ 1 5 1 ]
  //: joint g204 (w77) @(2376, 422) /w:[ 6 8 -1 5 ]
  OrMos g251 (.A(w237), .B(w91), .Z(w241));   //: @(2833, 466) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g97 (.A(w110), .B(w56), .Z(w137));   //: @(1193, 341) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: joint g120 (w69) @(1292, 356) /w:[ 2 4 -1 1 ]
  //: joint g66 (w48) @(785, 311) /w:[ 2 1 -1 4 ]
  OrMos g184 (.A(w149), .B(w74), .Z(w183));   //: @(2076, 350) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  //: joint g235 (w83) @(2617, 456) /w:[ 6 8 -1 5 ]
  //: joint g260 (w97) @(2975, 500) /w:[ 2 4 -1 1 ]
  OrMos g12 (.A(w132), .B(w61), .Z(w30));   //: @(418, 257) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g18 (w8) @(179, 228) /w:[ 2 4 -1 1 ]
  OrMos g226 (.A(w115), .B(w82), .Z(w223));   //: @(2539, 441) /symbol:3101448544 /sn:0 /w:[ 1 5 1 ]
  OrMos g283 (.A(w244), .B(w96), .Z(w181));   //: @(3130, 449) /symbol:3101448544 /sn:0 /w:[ 1 13 1 ]
  OrMos g108 (.A(w141), .B(w54), .Z(w52));   //: @(1032, 313) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g191 (.A(w180), .B(w80), .Z(w192));   //: @(2293, 435) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  //: joint g219 (w81) @(2436, 399) /w:[ 14 16 -1 13 ]
  OrMos g239 (.A(w228), .B(w84), .Z(w232));   //: @(2709, 456) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g134 (.A(w148), .B(w59), .Z(w115));   //: @(1472, 361) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g242 (.A(w226), .B(w84), .Z(w234));   //: @(2709, 400) /symbol:3101448544 /sn:0 /w:[ 1 13 0 ]
  //: joint g281 (w96) @(3089, 482) /w:[ 10 12 -1 9 ]
  //: OUT g4 (bin) @(3367,475) /sn:0 /w:[ 0 ]
  OrMos g154 (.A(w164), .B(w139), .Z(w167));   //: @(1746, 353) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g237 (.A(w220), .B(w93), .Z(w227));   //: @(2770, 475) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g58 (.A(w31), .B(w47), .Z(w88));   //: @(765, 259) /symbol:3101448544 /sn:0 /w:[ 0 0 0 ]
  OrMos g186 (.A(w174), .B(w72), .Z(w180));   //: @(2229, 430) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  //: joint g112 (w69) @(1292, 343) /w:[ 6 8 -1 5 ]
  OrMos g268 (.A(w243), .B(w95), .Z(w253));   //: @(2954, 420) /symbol:3101448544 /sn:0 /w:[ 0 17 1 ]
  //: joint g76 (w51) @(878, 321) /w:[ 1 2 -1 8 ]
  OrMos g211 (.A(w201), .B(w81), .Z(w204));   //: @(2477, 450) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g292 (.A(w198), .B(w41), .Z(w225));   //: @(3193, 482) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  //: joint g157 (w70) @(1847, 410) /w:[ 1 2 -1 8 ]
  OrMos g163 (.A(w169), .B(w193), .Z(w170));   //: @(1950, 410) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: joint g238 (w91) @(2792, 485) /w:[ 2 4 -1 1 ]
  OrMos g263 (.A(w245), .B(w95), .Z(w247));   //: @(2954, 448) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  //: joint g259 (w90) @(2853, 476) /w:[ 6 8 -1 5 ]
  //: joint g64 (w47) @(740, 306) /w:[ 6 5 -1 8 ]
  //: joint g166 (w75) @(1967, 420) /w:[ 2 4 -1 1 ]
  //: joint g294 (w41) @(3152, 501) /w:[ 6 8 -1 5 ]
  OrMos g274 (.A(w251), .B(w97), .Z(w257));   //: @(3003, 481) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g121 (.A(w142), .B(w69), .Z(w146));   //: @(1333, 351) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  OrMos g206 (.A(w199), .B(w79), .Z(w210));   //: @(2355, 370) /symbol:3101448544 /sn:0 /w:[ 0 13 1 ]
  //: joint g241 (w84) @(2668, 419) /w:[ 10 12 -1 9 ]
  OrMos g28 (.A(w13), .B(w7), .Z(w14));   //: @(174, 218) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g225 (.A(w207), .B(w83), .Z(w216));   //: @(2658, 465) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  //: joint g272 (w100) @(3027, 477) /w:[ 10 12 -1 9 ]
  OrMos g265 (.A(w246), .B(w95), .Z(w251));   //: @(2954, 476) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  OrMos g177 (.A(w143), .B(w75), .Z(w155));   //: @(2006, 387) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  //: joint g192 (w80) @(2252, 412) /w:[ 6 8 -1 5 ]
  OrMos g208 (.A(w114), .B(w77), .Z(w208));   //: @(2417, 403) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  OrMos g7 (.A(w16), .B(w3), .Z(w5));   //: @(257, 200) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  //: joint g262 (w90) @(2853, 448) /w:[ 10 12 -1 9 ]
  OrMos g149 (.A(w154), .B(w65), .Z(w161));   //: @(1688, 334) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  OrMos g286 (.A(w261), .B(w96), .Z(w176));   //: @(3130, 491) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  //: joint g207 (w79) @(2314, 403) /w:[ 10 12 -1 9 ]
  OrMos g296 (.A(w263), .B(w41), .Z(w248));   //: @(3193, 440) /symbol:3101448544 /sn:0 /w:[ 1 17 0 ]
  //: joint g48 (w40) @(590, 263) /w:[ 6 8 -1 5 ]
  //: joint g200 (w77) @(2376, 450) /w:[ 2 4 -1 1 ]
  //: joint g276 (w96) @(3089, 510) /w:[ 2 4 -1 1 ]
  OrMos g17 (.A(w21), .B(w42), .Z(w33));   //: @(477, 248) /symbol:3101448544 /sn:0 /w:[ 1 0 1 ]
  OrMos g29 (.A(w17), .B(w38), .Z(w20));   //: @(302, 247) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  //: joint g25 (w38) @(270, 252) /w:[ 2 4 -1 1 ]
  OrMos g271 (.A(w242), .B(w100), .Z(w249));   //: @(3068, 500) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g273 (.A(w215), .B(w97), .Z(w255));   //: @(3003, 467) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  OrMos g174 (.A(w178), .B(w193), .Z(w149));   //: @(1950, 340) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  OrMos g253 (.A(w222), .B(w90), .Z(w238));   //: @(2894, 429) /symbol:3101448544 /sn:0 /w:[ 1 13 1 ]
  OrMos g248 (.A(w229), .B(w90), .Z(w233));   //: @(2894, 485) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g80 (.A(w89), .B(w53), .Z(w107));   //: @(1086, 283) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  OrMos g94 (.A(w113), .B(w56), .Z(w127));   //: @(1193, 328) /symbol:3101448544 /sn:0 /w:[ 0 5 1 ]
  //: joint g193 (w72) @(2188, 379) /w:[ 10 12 -1 9 ]
  OrMos g202 (.A(w202), .B(w79), .Z(w206));   //: @(2355, 412) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  //: joint g270 (w100) @(3027, 505) /w:[ 2 4 -1 1 ]
  OrMos g21 (.A(w10), .B(w11), .Z(w43));   //: @(353, 224) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  OrMos g159 (.A(w167), .B(w68), .Z(w171));   //: @(1821, 358) /symbol:3101448544 /sn:0 /w:[ 1 5 1 ]
  OrMos g172 (.A(w159), .B(w74), .Z(w163));   //: @(2076, 420) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g232 (.A(w219), .B(w86), .Z(w226));   //: @(2598, 390) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  OrMos g256 (.A(w236), .B(w90), .Z(w245));   //: @(2894, 443) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  //: joint g41 (w156) @(513, 258) /w:[ 4 6 -1 3 ]
  //: joint g141 (w62) @(1523, 385) /w:[ 2 4 -1 1 ]
  //: joint g155 (w65) @(1647, 339) /w:[ 6 8 -1 5 ]
  //: joint g287 (w96) @(3089, 496) /w:[ 6 8 -1 5 ]
  OrMos g123 (.A(w147), .B(w69), .Z(w111));   //: @(1333, 295) /symbol:3101448544 /sn:0 /w:[ 0 13 1 ]
  OrMos g151 (.A(w153), .B(w139), .Z(w162));   //: @(1746, 395) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g90 (w55) @(1098, 328) /w:[ 6 8 -1 5 ]
  //: joint g222 (w86) @(2557, 465) /w:[ 2 4 -1 1 ]
  OrMos g82 (.A(w52), .B(w53), .Z(w108));   //: @(1084, 318) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  OrMos g128 (.A(w152), .B(w59), .Z(w57));   //: @(1472, 321) /symbol:3101448544 /sn:0 /w:[ 0 15 1 ]
  OrMos g243 (.A(w227), .B(w91), .Z(w229));   //: @(2833, 480) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  OrMos g33 (.A(w102), .B(w94), .Z(w130));   //: @(973, 321) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  OrMos g91 (.A(w107), .B(w56), .Z(w147));   //: @(1193, 290) /symbol:3101448544 /sn:0 /w:[ 1 11 1 ]
  //: joint g269 (w95) @(2913, 453) /w:[ 10 12 -1 9 ]
  OrMos g49 (.A(w36), .B(w40), .Z(w141));   //: @(625, 272) /symbol:3101448544 /sn:0 /w:[ 0 3 0 ]
  OrMos g137 (.A(w111), .B(w59), .Z(w158));   //: @(1472, 305) /symbol:3101448544 /sn:0 /w:[ 0 17 1 ]
  OrMos g198 (.A(w192), .B(w79), .Z(w197));   //: @(2355, 440) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g51 (.A(w78), .B(w50), .Z(w104));   //: @(859, 253) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g158 (.A(w66), .B(w70), .Z(w169));   //: @(1888, 405) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  OrMos g89 (.A(w103), .B(w55), .Z(w116));   //: @(1128, 299) /symbol:3101448544 /sn:0 /w:[ 1 9 1 ]
  //: joint g217 (w82) @(2498, 460) /w:[ 2 4 -1 1 ]
  OrMos g2 (.A(w9), .B(w6), .Z(w13));   //: @(132, 196) /symbol:3101448544 /sn:0 /w:[ 3 1 0 ]
  OrMos g77 (.A(w39), .B(w94), .Z(w134));   //: @(973, 293) /symbol:3101448544 /sn:0 /w:[ 0 5 1 ]
  OrMos g290 (.A(w181), .B(w41), .Z(w112));   //: @(3193, 454) /symbol:3101448544 /sn:0 /w:[ 0 15 0 ]
  //: joint g148 (w139) @(1705, 400) /w:[ 2 4 -1 1 ]
  OrMos g213 (.A(w205), .B(w81), .Z(w209));   //: @(2477, 394) /symbol:3101448544 /sn:0 /w:[ 0 15 1 ]
  //: joint g252 (w91) @(2792, 471) /w:[ 6 8 -1 5 ]
  OrMos g72 (.A(w71), .B(w51), .Z(w102));   //: @(910, 316) /symbol:3101448544 /sn:0 /w:[ 0 0 0 ]
  OrMos g203 (.A(w197), .B(w77), .Z(w201));   //: @(2417, 445) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g161 (.A(w161), .B(w70), .Z(w173));   //: @(1888, 349) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g182 (.A(w188), .B(w76), .Z(w177));   //: @(2138, 369) /symbol:3101448544 /sn:0 /w:[ 1 9 1 ]
  OrMos g196 (.A(w105), .B(w80), .Z(w200));   //: @(2293, 393) /symbol:3101448544 /sn:0 /w:[ 1 9 1 ]
  //: joint g152 (w68) @(1780, 405) /w:[ 1 2 -1 8 ]
  //: joint g189 (w80) @(2252, 440) /w:[ 2 4 -1 1 ]
  OrMos g246 (.A(w232), .B(w93), .Z(w237));   //: @(2770, 461) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  //: joint g255 (w91) @(2792, 443) /w:[ 10 12 -1 9 ]
  OrMos g288 (.A(w166), .B(w41), .Z(w191));   //: @(3193, 510) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g10 (.A(w14), .B(w8), .Z(w27));   //: @(216, 223) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g212 (w81) @(2436, 427) /w:[ 6 8 -1 5 ]
  OrMos g32 (.A(w30), .B(w42), .Z(w32));   //: @(477, 262) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  //: joint g27 (w11) @(323, 229) /w:[ 1 2 -1 4 ]
  //: joint g199 (w79) @(2314, 417) /w:[ 6 8 -1 5 ]
  //: joint g187 (w72) @(2188, 407) /w:[ 6 8 -1 5 ]
  //: joint g240 (w84) @(2668, 461) /w:[ 6 8 -1 5 ]
  OrMos g9 (.A(w0), .B(w38), .Z(w10));   //: @(304, 219) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g57 (.A(w46), .B(w47), .Z(w78));   //: @(765, 245) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g142 (.A(w60), .B(w62), .Z(w157));   //: @(1564, 380) /symbol:3101448544 /sn:0 /w:[ 1 3 1 ]
  OrMos g71 (.A(w101), .B(w51), .Z(w39));   //: @(910, 288) /symbol:3101448544 /sn:0 /w:[ 1 5 1 ]
  //: joint g295 (w41) @(3152, 459) /w:[ 14 16 -1 13 ]
  //: joint g145 (w65) @(1647, 395) /w:[ 2 4 -1 1 ]
  OrMos g73 (.A(w99), .B(w94), .Z(w103));   //: @(973, 277) /symbol:3101448544 /sn:0 /w:[ 1 9 0 ]
  OrMos g42 (.A(w32), .B(w156), .Z(w36));   //: @(548, 267) /symbol:3101448544 /sn:0 /w:[ 0 0 1 ]
  assign {w41, w96, w100, w97, w95, w90, w91, w93, w84, w83, w86, w82, w81, w77, w79, w80, w72, w76, w74, w75, w193, w70, w68, w139, w65, w63, w62, w60, w59, w58, w69, w133, w56, w55, w53, w54, w94, w51, w50, w48, w47, w67, w64, w19, w40, w156, w42, w61, w11, w38, w3, w18, w8, w7, w9, w6, w29, w28, w25, w22} = pos; //: CONCAT g1713  @(20,452) /sn:0 /R:2 /w:[ 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 13 9 9 0 0 5 0 0 0 13 0 0 13 0 0 0 13 9 9 5 9 0 5 1 0 9 9 0 9 0 0 0 0 0 0 0 0 0 0 1 1 ] /dr:0 /tp:0 /drp:0
  OrMos g180 (.A(w155), .B(w74), .Z(w179));   //: @(2076, 392) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  //: joint g74 (w51) @(878, 293) /w:[ 4 6 -1 3 ]
  OrMos g168 (.A(w175), .B(w193), .Z(w105));   //: @(1950, 368) /symbol:3101448544 /sn:0 /w:[ 0 5 0 ]
  //: joint g181 (w76) @(2097, 402) /w:[ 6 8 -1 5 ]
  //: joint g117 (w58) @(1367, 361) /w:[ 1 2 -1 12 ]
  //: joint g79 (w94) @(942, 282) /w:[ 8 10 -1 7 ]
  OrMos g194 (.A(w183), .B(w72), .Z(w199));   //: @(2229, 360) /symbol:3101448544 /sn:0 /w:[ 1 13 1 ]
  OrMos g215 (.A(w208), .B(w81), .Z(w213));   //: @(2477, 408) /symbol:3101448544 /sn:0 /w:[ 1 11 0 ]
  OrMos g36 (.A(w44), .B(w67), .Z(w85));   //: @(721, 296) /symbol:3101448544 /sn:0 /w:[ 0 3 1 ]
  OrMos g216 (.A(w211), .B(w81), .Z(w215));   //: @(2477, 422) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g125 (.A(w144), .B(w58), .Z(w150));   //: @(1408, 343) /symbol:3101448544 /sn:0 /w:[ 0 5 1 ]
  OrMos g144 (.A(w157), .B(w63), .Z(w160));   //: @(1628, 385) /symbol:3101448544 /sn:0 /w:[ 0 0 1 ]
  //: joint g178 (w76) @(2097, 430) /w:[ 2 4 -1 1 ]
  //: joint g81 (w94) @(942, 298) /w:[ 4 6 -1 3 ]
  //: joint g275 (w97) @(2975, 486) /w:[ 6 8 -1 5 ]
  //: joint g22 (w3) @(227, 247) /w:[ 2 4 -1 1 ]
  OrMos g45 (.A(w37), .B(w40), .Z(w73));   //: @(625, 244) /symbol:3101448544 /sn:0 /w:[ 0 11 0 ]
  OrMos g70 (.A(w88), .B(w51), .Z(w99));   //: @(910, 272) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  OrMos g282 (.A(w253), .B(w100), .Z(w263));   //: @(3068, 430) /symbol:3101448544 /sn:0 /w:[ 0 13 0 ]
  OrMos g114 (.A(w127), .B(w133), .Z(w140));   //: @(1264, 333) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  OrMos g209 (.A(w206), .B(w77), .Z(w211));   //: @(2417, 417) /symbol:3101448544 /sn:0 /w:[ 0 7 1 ]
  OrMos g279 (.A(w257), .B(w100), .Z(w261));   //: @(3068, 486) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  OrMos g229 (.A(w223), .B(w86), .Z(w224));   //: @(2598, 446) /symbol:3101448544 /sn:0 /w:[ 0 7 0 ]
  assign bin = {w191, w235, w225, w247, w112, w248}; //: CONCAT g30  @(3242,475) /sn:0 /w:[ 1 1 1 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  OrMos g164 (.A(w172), .B(w68), .Z(w178));   //: @(1821, 330) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  //: joint g289 (w41) @(3152, 487) /w:[ 10 12 -1 9 ]
  OrMos g118 (.A(w138), .B(w69), .Z(w135));   //: @(1331, 324) /symbol:3101448544 /sn:0 /w:[ 0 11 1 ]

endmodule
//: /netlistEnd

//: /hdlBegin signal
//: interface  /sz:(129, 107) /bd:[ Lo0<p2(48/107) Lo1<p1(32/107) Lo2<p(16/107) Ro0<clk(26/107) Ro1<fdbks(10/107) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls
module signal(p);
  output clk;     // this will provide a intermittent signal as clock (t)
  output p;       // this will provide the value of the s(t)
  output p1;      // this will be used for setting on boot time all the values 
  output p2;      // this will be used for setting on boot time the values 
  output fdbks;   // this will be zero on boot time 
  reg p;
  reg p1;
  reg p2;
  reg clk;
  reg fdbks;
  
  initial
    begin
      fdbks = 0; // setting all to zero 
      clk = 0;
      p = 0;
      p1 = 0;
      p2 = 0;
      
      $tkg$wait(500);
      repeat (58)
      begin
        #100 clk = !clk;  // Setting all the cirquit to zero.
        #100 clk = !clk;  // by shifting a zero value on the shift register.
      end
      $tkg$wait(200);
      p = 1;              // using p1 p2 p3 a single pulse of 1 is send to each shift register 
      #100 clk = !clk;    // of second minutes hours.
      #100 clk = !clk; 
      $tkg$wait(100);
      p = 0;    
      #100 clk = !clk;
      #100 clk = !clk;
      p1 = 1;
      p2 = 1;
      #100 clk = !clk;
      #100 clk = !clk;
      p1 = 0;
      p2 = 0;
      fdbks = 1;          // turning fdbks to zero ve comunicate that boot's time is done         
      forever
      begin              // This is the main signal, it will run  forever!  
        $tkg$wait(500);
        clk = !clk;
      end
    end

endmodule
//: /hdlEnd


`timescale 1ns/1ns

//: /netlistBegin D_FF
module D_FF(NQ, Q, CP, D);
//: interface  /sz:(40, 56) /bd:[ Li0>CP(37/56) Li1>D(13/56) Ro0<NQ(37/56) Ro1<Q(14/56) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(438,209)(390,209){1}
//: {2}(386,209)(376,209){3}
//: {4}(388,211)(388,236)(321,236)(321,256)(331,256){5}
output NQ;    //: /sn:0 {0}(438,270)(385,270){1}
//: {2}(383,268)(383,246)(319,246)(319,222)(334,222){3}
//: {4}(381,270)(373,270){5}
input D;    //: /sn:0 {0}(-143,236)(-109,236)(-109,195)(41,195){1}
input CP;    //: /sn:0 {0}(-139,296)(-108,296)(-108,330)(-93,330){1}
wire w6;    //: /sn:0 {0}(134,222)(114,222)(114,237)(204,237)(204,270)(176,270){1}
wire w15;    //: /sn:0 {0}(150,330)(214,330)(214,285){1}
//: {2}(216,283)(238,283){3}
//: {4}(214,281)(214,222)(238,222){5}
wire w1;    //: /sn:0 {0}(-22,330)(-8,330){1}
//: {2}(-4,330)(79,330){3}
//: {4}(-6,328)(-6,307)(-6,307)(-6,285){5}
//: {6}(-4,283)(41,283){7}
//: {8}(-6,281)(-6,222)(41,222){9}
wire w8;    //: /sn:0 {0}(134,256)(116,256)(116,243)(191,243)(191,211){1}
//: {2}(191,207)(191,195)(238,195){3}
//: {4}(189,209)(176,209){5}
wire w17;    //: /sn:0 {0}(238,256)(228,256)(228,243)(295,243)(295,211){1}
//: {2}(295,207)(295,195)(334,195){3}
//: {4}(293,209)(280,209){5}
wire w2;    //: /sn:0 {0}(41,256)(31,256)(31,243)(98,243)(98,211){1}
//: {2}(98,207)(98,195)(134,195){3}
//: {4}(96,209)(83,209){5}
wire w12;    //: /sn:0 {0}(331,283)(295,283)(295,270)(280,270){1}
wire w5;    //: /sn:0 {0}(83,270)(119,270)(119,283)(134,283){1}
//: enddecls

  //: OUT g4 (NQ) @(435,270) /sn:0 /w:[ 0 ]
  NotMos g8 (.A(CP), .Z(w1));   //: @(-92, 314) /sz:(69, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  //: OUT g3 (Q) @(435,209) /sn:0 /w:[ 0 ]
  NandMos g13 (.B(w15), .A(w17), .Z(w12));   //: @(239, 251) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>0 Ro0<1 ]
  //: IN g2 (CP) @(-141,296) /sn:0 /w:[ 0 ]
  //: IN g1 (D) @(-145,236) /sn:0 /w:[ 0 ]
  NandMos g11 (.B(w12), .A(Q), .Z(NQ));   //: @(332, 251) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>5 Ro0<5 ]
  //: joint g16 (w1) @(-6, 330) /w:[ 2 4 1 -1 ]
  NandMos g10 (.B(w5), .A(w8), .Z(w6));   //: @(135, 251) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 ]
  //: joint g19 (w8) @(191, 209) /w:[ -1 2 4 1 ]
  NandMos g6 (.B(w1), .A(D), .Z(w2));   //: @(42, 190) /sz:(40, 40) /sn:0 /p:[ Li0>9 Li1>1 Ro0<5 ]
  NandMos g7 (.B(w1), .A(w2), .Z(w5));   //: @(42, 251) /sz:(40, 40) /sn:0 /p:[ Li0>7 Li1>0 Ro0<0 ]
  NandMos g9 (.B(w6), .A(w2), .Z(w8));   //: @(135, 190) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>3 Ro0<5 ]
  NotMos g15 (.A(w1), .Z(w15));   //: @(80, 314) /sz:(69, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: joint g20 (w15) @(214, 283) /w:[ 2 4 -1 1 ]
  //: joint g17 (w1) @(-6, 283) /w:[ 6 8 -1 5 ]
  NandMos g14 (.B(NQ), .A(w17), .Z(Q));   //: @(335, 190) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>3 Ro0<3 ]
  //: joint g21 (w17) @(295, 209) /w:[ -1 2 4 1 ]
  //: joint g23 (NQ) @(383, 270) /w:[ 1 2 4 -1 ]
  //: joint g22 (Q) @(388, 209) /w:[ 1 -1 2 4 ]
  NandMos g12 (.B(w15), .A(w8), .Z(w17));   //: @(239, 190) /sz:(40, 40) /sn:0 /p:[ Li0>5 Li1>3 Ro0<5 ]
  //: joint g18 (w2) @(98, 209) /w:[ -1 2 4 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin AndMos
module AndMos(B, Z, A);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(187,223)(213,223)(213,223)(276,223){1}
//: {2}(278,221)(278,216)(293,216){3}
//: {4}(278,225)(278,228)(293,228){5}
input A;    //: /sn:0 {0}(179,173)(210,173){1}
output Z;    //: /sn:0 {0}(480,202)(522,202)(522,202)(537,202){1}
wire w3;    //: /sn:0 {0}(293,165)(278,165)(278,170){1}
//: {2}(276,172)(208,172){3}
//: {4}(278,174)(278,177)(293,177){5}
wire w2;    //: /sn:0 {0}(418,204)(370,204)(370,226)(355,226){1}
wire w5;    //: /sn:0 {0}(418,192)(370,192)(370,175)(355,175){1}
//: enddecls

  //: joint g4 (B) @(278, 223) /w:[ -1 2 1 4 ]
  //: joint g3 (w3) @(278, 172) /w:[ -1 1 2 4 ]
  NorMos g2 (.B(w2), .A(w5), .Z(Z));   //: @(419, 180) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  NorMos g1 (.B(w3), .A(w3), .Z(w5));   //: @(294, 153) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>5 Li1>0 Ro0<1 ]
  //: IN g6 (B) @(185,223) /sn:0 /w:[ 0 ]
  //: OUT g7 (Z) @(534,202) /sn:0 /w:[ 1 ]
  //: IN g5 (A) @(177,173) /sn:0 /w:[ 0 ]
  NorMos g0 (.B(B), .A(B), .Z(w2));   //: @(294, 204) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>5 Li1>3 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin NotMos
module NotMos(A, Z);
//: interface  /sz:(69, 40) /bd:[ Li0>A(16/40) Ro0<Z(16/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w4;    //: /sn:0 {0}(264,92)(264,132){1}
input A;    //: /sn:0 {0}(176,168)(240,168)(240,168)(241,168){1}
//: {2}(243,166)(243,140)(250,140){3}
//: {4}(243,170)(243,197)(250,197){5}
supply0 w111;    //: /sn:0 {0}(264,232)(264,206){1}
output Z;    //: /sn:0 {0}(264,149)(264,164){1}
//: {2}(266,166)(288,166)(288,166)(323,166){3}
//: {4}(264,168)(264,189){5}
//: enddecls

  _GGNMOS #(2, 1) g1978 (.Z(Z), .S(w111), .G(A));   //: @(258,197) /sn:0 /w:[ 5 1 5 ]
  _GGPMOS #(2, 1) g1979 (.Z(Z), .S(w4), .G(A));   //: @(258,140) /sn:0 /w:[ 0 1 3 ]
  //: IN g1 (A) @(174,168) /sn:0 /w:[ 0 ]
  //: joint g1980 (Z) @(264, 166) /w:[ 2 1 -1 4 ]
  //: VDD g1976 (w4) @(275,92) /sn:0 /w:[ 0 ]
  //: joint g1977 (A) @(243, 168) /w:[ -1 2 1 4 ]
  //: GROUND g1981 (w111) @(264,238) /sn:0 /w:[ 0 ]
  //: OUT g0 (Z) @(320,166) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin NandMos
module NandMos(B, Z, A);
//: interface  /sz:(40, 40) /bd:[ Li0>B(29/40) Li1>A(10/40) Ro0<Z(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(185,246)(262,246){1}
//: {2}(264,244)(264,239)(279,239){3}
//: {4}(264,248)(264,251)(279,251){5}
input A;    //: /sn:0 {0}(279,188)(264,188)(264,193){1}
//: {2}(262,195)(185,195){3}
//: {4}(264,197)(264,200)(279,200){5}
output Z;    //: /sn:0 {0}(564,225)(625,225)(625,224)(636,224){1}
wire w0;    //: /sn:0 {0}(493,225)(466,225){1}
wire w2;    //: /sn:0 {0}(404,227)(356,227)(356,249)(341,249){1}
wire w5;    //: /sn:0 {0}(404,215)(356,215)(356,198)(341,198){1}
//: enddecls

  NotMos g8 (.A(w0), .Z(Z));   //: @(494, 209) /sz:(69, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: joint g4 (B) @(264, 246) /w:[ -1 2 1 4 ]
  //: joint g3 (A) @(264, 195) /w:[ -1 1 2 4 ]
  NorMos g2 (.B(w2), .A(w5), .Z(w0));   //: @(405, 203) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  NorMos g1 (.B(A), .A(A), .Z(w5));   //: @(280, 176) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>5 Li1>0 Ro0<1 ]
  //: IN g6 (B) @(183,246) /sn:0 /w:[ 0 ]
  //: OUT g7 (Z) @(633,224) /sn:0 /w:[ 1 ]
  //: IN g5 (A) @(183,195) /sn:0 /w:[ 3 ]
  NorMos g0 (.B(B), .A(B), .Z(w2));   //: @(280, 227) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>5 Li1>3 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin PosBin12
module PosBin12(bin, pos);
//: interface  /sz:(100, 40) /bd:[ Li0>pos[11:0](16/40) Ro0<bin[3:0](16/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [3:0] bin;    //: /sn:0 {0}(#:765,316)(830,316){1}
input [11:0] pos;    //: /sn:0 {0}(#:74,332)(#:106,332){1}
wire w6;    //: /sn:0 {0}(307,337)(293,337)(293,337)(270,337){1}
//: {2}(268,335)(268,312)(304,312){3}
//: {4}(266,337)(135,337)(135,337)(112,337){5}
wire w7;    //: /sn:0 {0}(112,357)(234,357)(234,357)(444,357){1}
wire w16;    //: /sn:0 {0}(417,283)(423,283)(423,282)(452,282){1}
wire w14;    //: /sn:0 {0}(337,332)(350,332)(350,337)(387,337){1}
wire w4;    //: /sn:0 {0}(202,302)(304,302){1}
wire w19;    //: /sn:0 {0}(660,372)(702,372)(702,331)(759,331){1}
wire w15;    //: /sn:0 {0}(334,307)(340,307)(340,302)(387,302){1}
wire w3;    //: /sn:0 {0}(112,367)(356,367)(356,367)(426,367){1}
//: {2}(430,367)(444,367){3}
//: {4}(428,365)(428,292)(452,292){5}
wire w0;    //: /sn:0 {0}(542,372)(532,372)(532,377)(522,377){1}
//: {2}(520,375)(520,317)(540,317){3}
//: {4}(518,377)(112,377){5}
wire w21;    //: /sn:0 {0}(482,287)(576,287)(576,296)(600,296){1}
wire w28;    //: /sn:0 {0}(112,317)(252,317){1}
wire w24;    //: /sn:0 {0}(642,317)(686,317)(686,311)(759,311){1}
wire w20;    //: /sn:0 {0}(417,342)(693,342)(693,321)(759,321){1}
wire w1;    //: /sn:0 {0}(119,277)(112,277){1}
wire w25;    //: /sn:0 {0}(282,322)(297,322)(297,327)(307,327){1}
wire w8;    //: /sn:0 {0}(387,347)(368,347)(368,347)(364,347){1}
//: {2}(362,345)(362,314){3}
//: {4}(364,312)(377,312)(377,312)(387,312){5}
//: {6}(362,310)(362,288)(387,288){7}
//: {8}(360,347)(112,347){9}
wire w30;    //: /sn:0 {0}(112,287)(138,287)(138,268)(172,268){1}
wire w22;    //: /sn:0 {0}(570,312)(612,312){1}
wire w17;    //: /sn:0 {0}(417,307)(488,307)(488,307)(540,307){1}
wire w12;    //: /sn:0 {0}(282,278)(315,278)(315,278)(387,278){1}
wire w2;    //: /sn:0 {0}(202,273)(210,273)(210,273)(252,273){1}
wire w11;    //: /sn:0 {0}(630,377)(610,377)(610,377)(579,377){1}
//: {2}(577,375)(577,360)(577,360)(577,324){3}
//: {4}(579,322)(612,322){5}
//: {6}(577,320)(577,306)(600,306){7}
//: {8}(577,379)(577,387)(112,387){9}
wire w10;    //: /sn:0 {0}(759,301)(710,301)(710,301)(630,301){1}
wire w13;    //: /sn:0 {0}(474,362)(527,362)(527,362)(542,362){1}
wire w27;    //: /sn:0 {0}(572,367)(619,367)(619,367)(630,367){1}
wire w29;    //: /sn:0 {0}(172,307)(158,307)(158,307)(150,307){1}
//: {2}(148,305)(148,278)(172,278){3}
//: {4}(146,307)(112,307){5}
wire w9;    //: /sn:0 {0}(252,327)(238,327){1}
//: {2}(236,325)(236,283)(252,283){3}
//: {4}(234,327)(130,327)(130,327)(112,327){5}
wire w26;    //: /sn:0 {0}(112,297)(157,297)(157,297)(172,297){1}
//: enddecls

  OrMos g8 (.A(w28), .B(w9), .Z(w25));   //: @(268, 322) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: OUT g4 (bin) @(827,316) /sn:0 /w:[ 1 ]
  //: joint g13 (w9) @(236, 327) /w:[ 1 2 4 -1 ]
  OrMos g3 (.A(w2), .B(w9), .Z(w12));   //: @(268, 278) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  //: joint g2 (w29) @(148, 307) /w:[ 1 2 4 -1 ]
  OrMos g1 (.A(w26), .B(w29), .Z(w4));   //: @(188, 302) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  OrMos g16 (.A(w16), .B(w3), .Z(w21));   //: @(468, 287) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g11 (.A(w15), .B(w8), .Z(w17));   //: @(403, 307) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  //: joint g28 (w0) @(520, 377) /w:[ 1 2 4 -1 ]
  OrMos g10 (.A(w12), .B(w8), .Z(w16));   //: @(403, 283) /symbol:3101448544 /sn:0 /w:[ 1 7 0 ]
  OrMos g19 (.A(w7), .B(w3), .Z(w13));   //: @(460, 362) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g27 (.A(w30), .B(w29), .Z(w2));   //: @(188, 273) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  assign {w11, w0, w3, w7, w8, w6, w9, w28, w29, w26, w30, w1} = pos; //: CONCAT g6  @(107,332) /sn:0 /R:2 /w:[ 9 5 0 0 9 5 5 0 5 0 0 1 1 ] /dr:0 /tp:1 /drp:0
  OrMos g9 (.A(w25), .B(w6), .Z(w14));   //: @(323, 332) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  OrMos g7 (.A(w4), .B(w6), .Z(w15));   //: @(320, 307) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]
  OrMos g20 (.A(w21), .B(w11), .Z(w10));   //: @(616, 301) /symbol:3101448544 /sn:0 /w:[ 1 7 1 ]
  OrMos g15 (.A(w14), .B(w8), .Z(w20));   //: @(403, 342) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: joint g31 (w8) @(362, 312) /w:[ 4 6 -1 3 ]
  //: joint g17 (w11) @(577, 377) /w:[ 1 2 -1 8 ]
  assign bin = {w19, w20, w24, w10}; //: CONCAT g25  @(764,316) /sn:0 /w:[ 0 1 1 1 0 ] /dr:1 /tp:1 /drp:1
  //: IN g5 (pos) @(72,332) /sn:0 /w:[ 0 ]
  //: joint g21 (w11) @(577, 322) /w:[ 4 6 -1 3 ]
  OrMos g24 (.A(w22), .B(w11), .Z(w24));   //: @(628, 317) /symbol:3101448544 /sn:0 /w:[ 1 5 0 ]
  OrMos g23 (.A(w13), .B(w0), .Z(w27));   //: @(558, 367) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: joint g22 (w3) @(428, 367) /w:[ 2 4 1 -1 ]
  OrMos g26 (.A(w27), .B(w11), .Z(w19));   //: @(646, 372) /symbol:3101448544 /sn:0 /w:[ 1 0 0 ]
  //: comment g0 @(363,415) /sn:0
  //: /line:"dec| bin  | Pos"
  //: /line:""
  //: /line:"00 | 0000 | 100000000000"
  //: /line:"01 | 0001 | 010000000000"
  //: /line:"02 | 0010 | 001000000000"
  //: /line:"03 | 0011 | 000100000000"
  //: /line:"04 | 0100 | 000010000000"
  //: /line:"05 | 0101 | 000001000000"
  //: /line:"06 | 0110 | 000000100000"
  //: /line:"08 | 1000 | 000000010000"
  //: /line:"09 | 1001 | 000000001000"
  //: /line:"10 | 1010 | 000000000100"
  //: /line:"11 | 1011 | 000000000010"
  //: /line:"12 | 1100 | 000000000001"
  //: /line:""
  //: /line:""
  //: /line:"13 | 1101"
  //: /line:"14 | 1110"
  //: /line:"15 | 1111"
  //: /line:""
  //: /end
  //: joint g12 (w8) @(362, 347) /w:[ 1 2 8 -1 ]
  //: joint g33 (w6) @(268, 337) /w:[ 1 2 4 -1 ]
  OrMos g30 (.A(w17), .B(w0), .Z(w22));   //: @(556, 312) /symbol:3101448544 /sn:0 /w:[ 1 3 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin OrMos
module OrMos(B, A, Z);
//: /symbol:3101448544
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(278,257)(406,257)(406,227)(430,227){1}
input A;    //: /sn:0 {0}(430,215)(408,215)(408,189)(278,189){1}
output Z;    //: /sn:0 {0}(621,225)(669,225){1}
wire w0;    //: /sn:0 {0}(550,225)(492,225){1}
//: enddecls

  //: IN g2 (B) @(276,257) /sn:0 /w:[ 0 ]
  NorMos g1998 (.B(B), .A(A), .Z(w0));   //: @(431, 203) /sz:(60, 40) /R:2 /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 ]
  //: IN g1 (A) @(276,189) /sn:0 /w:[ 1 ]
  NotMos g2004 (.A(w0), .Z(Z));   //: @(551, 209) /sz:(69, 40) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: OUT g0 (Z) @(666,225) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

